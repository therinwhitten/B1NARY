    ����          =B1NARY, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   B1NARY.DataPersistence.SaveSlot   datascriptPositionimagefileInfo+SerializableSlot+<LastSaved>k__BackingField*SerializableSlot+<TimeUsed>k__BackingFieldSerializableSlot+fileInfo  $B1NARY.DataPersistence.SaveSlot+Data   .B1NARY.DataPersistence.SaveSlot+ScriptPosition   System.IO.FileInfoSystem.IO.FileInfo   	   	   	   	   I��~�ڈ2��    	      $B1NARY.DataPersistence.SaveSlot+Data   choicestringsboolsintsfloats�System.Collections.Generic.Dictionary`2[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[B1NARY.Scripting.ScriptLine, B1NARY, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]�System.Collections.Generic.Dictionary`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]�System.Collections.Generic.Dictionary`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.Boolean, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]�System.Collections.Generic.Dictionary`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]�System.Collections.Generic.Dictionary`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.Single, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   	   	   		   	
   	      .B1NARY.DataPersistence.SaveSlot+ScriptPosition   	sceneNamedocumentPathlastLineSystem.IO.FileInfoB1NARY.Scripting.ScriptLine         Times Square	   ����B1NARY.Scripting.ScriptLine   lineDataIndextype  B1NARY.Scripting.ScriptLine+Type         SNew York City in Times Square: the year is 2040. Midday on a blistering Summer Day.   ���� B1NARY.Scripting.ScriptLine+Type   value__           �� �PNG

   IHDR     U   ��W#   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^佅Y�����o�35�U���T�L�233333�l������̶%ْm�bx����H�TruU���NM��TD�232#��|'ND����_�+������������������������������w��o?�g�
�>���߬Ś9��c�y�`�s��a}$wO���rBo5 ¶���Hs�@��cd������F��s��L�����A�w�"ǧ��������3h!�g���;�|�~�sڃ<�礛<En@����grI6��g�4��=6?!ϐ���ϑ�3��H>�e��O���q=Ȋ�US����׊�w��g��#;a�)r��]��K�w����DA�	ޗ�����q��qe�Y@I��8J�������<�<�( *��"mjF�.jJH�(jˀ�
��rU�h�ES�0�kF�R;��-�#h�%�����oƃ��5���A[��t�h<lչ�b:���P����~������M\��~n~'�i\��QT��,���=(�z ���=EI�u�(������|A ��u������ҌL�zd�U#�V)��"�BbO� �H,"F"ro�w� t{ B� t�?�H�f?�ma����m|���->��������[灰��]㎐5�Y偐��_��e�],D�pE�J7D�rG�j¿�Z����kl�@�VOn���nx����8
�������Xl����X���T���t8l�D��l$n���Ѱ����p��K��}!��$�Ϗ�`{&���׋���H�:a��<��!���!�:��qȟpz0x���� \��K|W�z�����}2�q�o7��P(���E�qy�G��dN���t�M���$�]L��tx]̀��,��́��\X�!Į����r�D�Kb�j�uH�j@�w���؄��dFp]��@nB'
�4��3�P�3�ʼQTs;�m��|Tmw��@3��nWi�%S���Zn5PS��\^K�iy]�Or�Md�n�lR�.$�$�	lK�4�bؾD��0r��l{BP��'h����9/S�]�?F��,�B�nOl���<�}}�	d��Z�s��I.my7RCIx7�Þ !�q������F�T�ۭN�鰱���+�8z�.����aŲC�;}+�~���5�a���o�M�?��?���_�_�ߗ������?_Ǜ��.�~�����������M�'��o�[�-����W�8�n���2�|!�����iHvnE��#d��	����� �G��X��-��m��* �" \�	� #������� �%�EPm M�+��HI@��8m���L!6D" ����aJ�����FX$���G ZuhfC��F���]��&eUIè�DyL?J�zQً����(�)���1��v�(�S���(�ec-�Jpj@���Y�!��x1	g�s<1Gb-�/�C�3�ۃ�-��N	���P�p:���!2����0J@�H�zJ E d�'��p�p(aDB�@��" |n�.j����O�所^��!8<& 2=�G ��7��������p�
~ۣ\���Ng�U�;�K��d�_J���4x�������_�?Ȧ ���Z�;U Ƶ��	��*��}���Hap�3�3��!+�9񏐟��)OQ�у��T����e`�2���_��a/�?��$ �*��l*�ɿ� H�OF!��
|f	_��z�g��� #�)��?� <� <z� X[���e?9�={ob�ƳX�� `�|���9�:���������~��_��W��/~����wx�^�k����W�_�+������W�������x��7��?�0S�[��_�����0���x��ӱ�뭈�S�T�6�=��?�
~�j��& ��
D���g�0����[����������HIQ+�&f����H �c�8�(����E &�L& U�`(	�D@KO e���M� hR����8�8ݫQ�o�B����ڥ'���~�f
K3�AI ����T���*y�=���Q�j+��oW�vyTJYq�ހ�.�BJ@!%���!� ׭Yw�i_�4�r��(B��\$^�D��ĝ��E��hD�P"�'��C�+Q;��#��� �B�NyL�)�v
�6
�@d l�`#ß"�j>X��I�*-��תĮ�D"r%b�'��x������ �RI��`ClO���tn��ĝ����E��<����Kqp��؟�����c,�1�m�6}k	��1�u,Vǂ_  ��q\?H��^���7�?�"8�|�;'"�1�8�~C?	���R����Z:��g0���o��@��mBn"̾Qw+�Ո�`�{���iP$�6!ſ�A�Hf�~YQml+�>1��R�Q�.����Bu�0j��Ip7p�2�_�]�p���=��@d[�7m[�k��J)�׬�6Q���@ۅJ��i��Hc[@	(��QJ��� ������ ���`�g��d;�M�y�M��?��`
�?5�	�û�ց��6Dߣ 4�	�C:���p��/s��ױ~�i,[�s�m·/�'o��{���	�?��?�W��~��_����W��o~�~�Ͽ����
^��k���?��w^����=���������o��)�{�+������W?���o��1�}�+Xqi������ #Y�, �T$���=� ��0�d�HO@~ E��f~� dpJ31NL�o���0C Ң�<C�,
��Y ��͢���c��Ч�I�W�o0Q�����q�b�M����`�  �@� 6z�O&" �`� �I���E���F���8�D��p�SM �v�ioQ���:j�Q�(ß��v	�P3�Vy��4�6��=�ܔ�j���2y�I��ҩL�(��U�߽�BX��(��H�. >��s��l�&d:�!Ͷ)7��|-I���x>	g�{�p<�G�u(
Q#s 1���a���h��SE�"j��(
��Hގ���ݔ����Dl�Ce t�7B6yQ����(}�Z��u^�^����F�FoDm�B�/���wx#p�7�w{�{���n� �a���-��H0�TH���`��WP �P �G���_��9o��WB`̟�<�~�3|����f��f��2����PXS ��9��7���qp��Ƙ�ڗ�7����>{~'~���KI
�+)
�ki�ߛ�����E�mo�#ؾ�N%�p.C�{�j�[�? �?����l{�#3�D>@vt���%�X���/�@e��
���IO�'���W���}�q
�Y ��v���/�e�H��;��Z�ſ��A5�*��'@�. �	@��4�]�?��ζ�P����A?�Y��f1�s�X�j�m(�����!�M�B�v���{B#-\�)��H�x���Ą�� G�4ܺ�s}( �kX��$�,ڋ�S7������gQ �������/��B���^��|��o^�%^����_�������ꗘ��Z�{�|���9Dc��G��˓X��~|���G�˟����,��c|��<��KF�W'ß?�;��'��K��ԟ+���""}�x�B0w��(bPOe@�S����	 �H��c/�Lf���0�I@��4_] &�L.����z��M����J�	�  �`�z�� � X$�U�4.Ra��e`\�!l�$���H��# �̴3�� H@����2�8��aJ )A��;��Y��V���*�HA�iU�*("�1=(��V��)�
�c=��T!պ�7�r-I���p1�ܖbO'"�d<���"�hb
A�ar(R�&�:�C)x�)
�C4�R�P
v"|��w�"|�¶y#|�7"�-��ԉ�꧈�@����wR"���{���~?V�>RV��G�m����P·��8C�A)ay��o��:��m�.+|��QJ���HqA`�/�ӥ{]�م;'(ǣT׻t��	W��V�-�^�1xߡc��,�����j�@���x(�ԖÉBb��7��KW����~��h����e_�}1�K�\��*D{0�}��J?%�C�>+�6�X;�\�Q�ȍ}���N��/�_�F����v)��\�m�0�%�����r=�@�𗐗����7eYM'	� �o"��R���֗����s-�������o��/����^��-��B^�� H��I����" Ya,�B�+�,����~	���N
@'��. m�
@=�+��Z �Tܼ���q�=v�u�Na��}���F|��R|���x�wS4��	�����|�_���2����������6l�v'Wy�jO+�Z��<���NdV�6+���0��x�����?�������x����F��ց,= ǃ���C ���(�cJX�P/�)���XH|��T��D��k��	�!��m�L�̸~% c`f��X0$`� d��a	Ȧ��̏� � �;�Hע� ]�� ���86@@��\ ��>�׬cY3��Jmw@?c3?{#��^oEjs���"��mR%ՐH@|���2��;�0�s� 4#�n2j�nW��Rd�*B��<$_�B�t$�OE��$�Q�G �2"q�c{�2@��D!�p$b��GP�C!�9�h��}�� D1ȣ��
%��9A��8��A���FA��`�F	<�#!�f�1��w`�;���3+t��Q��7�z1�Us����.���|1N�<���_]��f!�6���(%�h�z(�C-�� �?��M�o��	~C^dY\/�[��ؿo��7�_��K���.F�C"�#ܵQ5��c�߈��V��<@Fx2��ω�B^��w�0����/f��/��Cy� �1�?��:
����(7r=n�� �.���(�7�����_�Vq���<����4ȶZ<���Zn�5��U�_����*��>H�'�2���P�-�|�0Qƅ~���� �o��`f�~-�Yd
z�g���U��
���Ax@hFX@�*���;)�q#g�{��{��ukמ��{�ݷ��K�!�� H����
�o�/��������ά��eѰ��gU�(
���6!ýՉ�� �)��	âv����_}�"���Ç��)��������ɍ!K���A�'�_�b5�i6�9�-/�N�7�hc0��/W"�`!�Ї����0|��"2	Y�"�|:����t�Fy҃�r�n�
��M��԰.��i��I�z�$@PMd���X~6K� ���d�"'~�P�Hn�7y����~V����/����-�m��1V�l���S ��)�1_�^ c<��ꔳa�DH�� �R���@z��Z�V�Ѳ�������{�I��;�5P�Q��C	} Chk�r_v5����9Z((M�������\�6�\�z.g=����Cƪ�!J� �(k��=�)�����;(�m�.Z���*�n=2�j��P��;���r��*F�|$_��{�!��S�p!�R��sI�?�@)�C��hD��|!�x�Q�9FY8AaGԡ0�(V�0��!r?ŀS!�@0�!��B$�G�w,�����#��$��~�ǩ0����������ҝ!���`��3�ݯ0�/'-�=�$��j2+�x\M"�j�����)A�H)� #�)�8���,��gb�t:����@�?A�)a���h��bGl�,
.��P���Qf���Q��ݦ�؟��#����DZ�)-�\~�+�����U�o[�`	�;�w(E�S9����Z�XV�	�H�mB*�~���T�1���#?����E)�(a�fR(�{Q�ۏ�<V�CܖX�s۩�`Pˑ5�&����\�ǂ߀��nK��� p�������Q�O��u��۷Z�Et�Ev�ʿB���_��2�Kb���(�퇱��P 6�"
@q(!�B���X�˼�<f��6:�m�j�) 9��s��$'�R ��moFD�JTZ�#�D�#1��#�!:���5��.��k.�$����;�C�nc��+X���߃_�Ǘ�/���w^�w� ��Ƀ�?
/�7��-�|�3�ZtgV���X\]�����*���b�5��� Db�;��+��߿G���������i� 7�n����_��l/m `�א�<o��~H b�8S�k��{�7�� ;�2b"+�"��_ ��Z��DRC��Jۤh�I�� DR ���1�1N b��b�}Q r) f��])8/@�<�~���?�����M $��c^	�>`"*�'P�P��?Q�c@� iȆ)���,�$��(ha�c���ި��>C:���ި�	�v	hܓ���T�ш�mb#)ݣ\���\
@�*���%��$���`7�C��n>D���z�C����P�,J@�c2�T!]$���7�*�׳I�"�$\�@��4�]LBܹx�2���E#�l�����bO�R����c(Ѭ���S�Q�H�_�/��q��X��w�����g��3�Y�Ɲ��{G"�t������x�ϙx1�=����Kq���I��E<o�������Z|�%�9)�ޔ �+�� J (nb�z>�+q�p�w�r.�g~λ��N��-8�.
�d8�q8�|F{����o���K���t�o��V6?A6�+��;%jp_�c"Y�G�T���2�?Iٟ�Ϫ?�>�Y��ڗJ??���-��tV�*�{�}�~�� �#	~�7��A����~�\?I����0C ����M\�e�6��u\�k
��J�� ����7��� 0��$���@	��Pd� �P�	�& �A>�_�m�?/x��4�R �( B��@�H �t�v��LC �) 1�h����jFTX=B����[
��߉� ��Y7
�-�m��U��a��]���:|��bM ^�Y	����_���_�^{�|��|l�{�W��ʪ\[����<_��3e�;Y�*�>�C�o��] >�;�~�s;\��ډL�H����ߋ\ڠ`�� ��r����f؛���`������@j��1�Hf��ҩ$ ���&�`�0A�����~g�;�O5D
,��#7�� 
������q�n��D�" ��@����A9C*e�����1$@Q:B��ԗ��EG�H ԡ��Q R�K�w��'�Q2�Ϗ��&c��Z"|m��>�2�����$=�R-��kY��J�0�A6�� ��E����G��kC��}丷P���R�l�@��ZdS��7�v2mK�nS�T�|��H!I���Hd %\IF<+�x�b�.�N��$\HTȼ�ās,�Y�x����e��Iس��O`�'�DV��D�o"C8���m$�6��������w9~��IIB��Z�"�&�_�kN��X5�!�f*��
N��~_�����r%^����e��(�
�r���q��@n��J X�O��9>�ߝ�%y?J��TJK:|o1�2���h���>���j_��/B����/SD;K�W(bܪ�^��E�OR���؂�`Xr""?���ũ=��P�3���Tp�(�3�e���$��� b,�c�-p]lnf�j��uߠ�<��@v�ꟕ���zM����gٵ �t��u��'�?:# ڮ �1�G���|V���l�B٦#�#����g���QO���P b&���*�����%wn���� �=㊃m�u�%�\y���Ĵ/���w��?��;����% ���e���?�����3|��X���[�K+�qu�'3[�QЍBqqe,έ	Â�w��}���!���Gx��S >Ùmw�x���!\��_! � �a>�|�L�?��d� �1�uR���]Hxl!��/$� H/ ��Q�Oƍ	0I�O�����8
@<C=�L"7�$b0� a20��-	0$�"�$ �nb�� HW�H�d `���I�R�3�e�'Q��pҦ�}O;F�Luڵ�����RF4��PB��Jh�FO��o+`�2��Vˬu���
(��Aq�SR��ە �z�p�� �7 ׭9�u�q�ܭ�T#ӡ�eH�SL�i���*3�*�7)��(�H�.�ZH��L�%		�
 �L���D�%�A{)��x��܎��z�1���"��.����U�O`Ǔh�}$���j>�fBn��٦#�.�w�a��p�l��Pb���;٬�3��[�#���������"\� �.��%~|?�S|�o�m���x��{]�~W���o�!��/Az�A�Ƞw*D��޵Qn��v����u�B���7F�W-�8�S��:$�7��`���c�� ���g8�?Fqr7J�d4?�Y��K�6F�� +]�r�,�W��^��8���i��?������\�8�\���lO�m�{���v�z����Q�e������ ȉ�) ����8?� (L0�'� � c�>�J�ۤ0�6?�Ou�O�o���Y�O, ��#���@�Q`M8�+cޜ���*
�|����x�7_���7/�/���X7� }�������|cvϲš���
�#�8�؝�ݰ�=f��o0���(�߿�w_�'6�#��=$�w"ӹ���ڀ@S�����
�y���d���	���c��h���a�g����F��S��<A�|)>]H�}�$?�=E���P�X�#����B9PǢ>�H��z̌;*�G� ��k��� ��DZt��dޞ��'J��wp�<(�$F��E�����nJ���L��L�PS��h����.�100$� �A� @����Rի��;�Q<{8�g�F�str��n%#J)�������Ȕ��QEI#��&cd|�4�U�J~�2�8���N
䌀�^�G�W3��f�yr�ވ\W�G ǥ��5ȼK	p*G��RE�S	R�"�.I�B�NI�V�I�d�5M�I1`p&���gx�3��ޟ�j<�a��<���&���=�W�GHP!�z��nC5��p�2����4�D�5��Rm���;�v�D�S.���R�x�BđX#S�"�8"�1��N��0p̄��3sY,py���~� ~����ې�@.kЭ
����6 \O��!�,���1Ԇ��v."�Y���/c�W λ�a^�0�ePg!%��}P��HiB*ImFfx+�>�b���P�؅R9�O�3�g��*w 5�0>��2 OD��������8b�Ч��� tp;��TU��T�Yo�7K�d��ȶ�w�7��ob�7c[���a��/���B��!�� J@QĠ�����ȏ!l�����M��#( �=��'!��wß��i��c!3�KMSb:�4a�! ��bq�J N�r���Vؼ�<�/?����a��������) ����k��~�+�����y7qv�'vwo��9��/��+3��k�����?LǗ�-��.�'������x��w�������:7��u���kA�]R:��ҥ|� �x2�t�2���H�d�����×����=F�7W^\yH�WRuR<��I������>�Ƒ�ۉ� "@��+�����d��%`bo�d2�c:*@�
L�`F� ~w�Pr�x{R�`�" `��D0��C2,��� �	�E�� 9��O i��  9���������C��F��d}O�B���ǣ|���(�j=��G�}D�m�2��le��2��0�Fm�Ӯ��p9����F�����>F��ۮ$ ק��.�&w�֤��pZ��v�D:E š�"��T�]6��ɷ�y_��&2Hm2��0M`JH'r�b��4V㩶k
��M�ߤ)���\�d$34��I�D���L�$�-�/�5���:�[���O���u�B�S6�]r�̠O�x� է�]�d�$�^�H�,C�[1���#�>��G����A	�"��H��A�L�>
P8�)����b��P�9���=�<?s�.���"���J?��~�?�O�����HkBfD����so{N�Ent����6d����ű��j_N����ϸ���*����\oF��0����ܗC�X��o�:6�@'��h���<���i�Ϡ�' z�K������hٞ��Az���	��T�\�����ꇾ�4(���@�d��2�5�1��T��Mc��F��^�J���*	��؇/ ���9v�1�r���r˖Y���g� ��,|祟� ������W~���˛���k�pa�7^�3��Ƿ1��EX��>,��V|q�?ݏ�����/v��g�/��NxG� �M���_��f{�ܬA��}6���؁4��pc�y�� � P
<ΓO���=F.�o��+�$d�>'���t#ˋv詑���dypE�)*��x�������C$�DH�;�юxO�{=D�oS(	~�
�H@ C?H�PB�,����<GWbѼ-�BիK �ބ�69ȉc��[�y	#ȥ�$�1��D>����4Fn�x	�sO��7 C����X�ͻ�GǇ�.F�@�.�z�����% ���xVCR�?d��*��	�c��_����=c��(�GI =���"�#xJ?A��tv�h=m�êQ!i��k�rȡ�" U� �_PJ�+���wP�P�w_��>���Z4�h���}B�"׳��Jҝ�(��Heh�9
y�/iyH���0�B�� �>њ�n���B�c�#�����52�����,5�b�N�����̠LdE/�� ��n�l������e��8e��2�S��Y<��[�,�
dT ;�Y$3��T�v�k��[�m��wX��A��@,�>�@n�󸜱�.sG��B��'�#�j���c9���#���&�RV��^�-�~�F䄵� �
�����](!�):2�P/Iy�(MCݧ~�)����P�7���!40�%|e7�T���t��v�y�=N������v�g;׻v�\�e�M��:?fP�� ����n0���=[�r����/U���mTN�-�_#���GT��T(7I��'�(z�&
�M��Q�� ��}ڇ���d�6R �z���NE���w�. Ѹ|�'O�ž}��i�9,]z�gR �: o��}u����j�K�%%��_��]����_�a��_���_�n�Q\]��˂qyU..�¥������l�[�{}�-�����Ϋ�b�'sp|����"�F#��	� ɑ?�w��'D�u�E@�C������a�������!�i�_B^�;������$խ]���`���!O�8s���q�Ľ]K���TD���"ІDVw�����
�t"I�2�7����i����r;�+�AW��C9�a�ǌ�� �Z��o@~���#�
��������/E�_vȑ ڮ ���1�H9�
�L�v%3Ul\��J�'�2@�vh�J�7Tȑl$����ʪ[�����T3lԤ��`�?b��Ɇ��#
 ����%��З��F���I�F�0����[�󧔀'�x�x��;�$���(>�i B��UO��ȲS�D �b( rb �`Q�C% E�c�=P ��M�E�w#
}��4ϳV�d��!ݹi�T�<N��°%鬤Sr( � �3:����2��)� iw)���ټ?����r[{,�2���!�&���H�|2�|�-��T0����TG��k>�9>��e��� ?�VQ^�*��\�hkd3�S����_�$�5���	|�D��)I�x$��J����M��2�r�dJD
eH����Hr*@��B���S�����(E�;����CA񯦨�#7���Q��I](K�F�^�W���*���ud^�:��B-�7F?��M�#hf跔�үЎ�W�/��p~����:%r)�WG����VP>I'����\���d���?�	~�16�]Q'��{�a�r��nc-��g��&���u���t-��n��1���Sc'��?���D�	�b�������H-����E����
"9Q��%Œ^���p�6?^#-��%� �� �<@BT+�B�P���n&lm48q�{���ƍg�t�̞�S>^��ߘ�?���g5p� ����Ӭ��˟�W�Ǧi�pc]
�m
ą����&7���fs,�~���>�x����{x�Oa�7�qp�Mx_*D��Z�ݨG�M+�n�wd:?�H��Y �Q2��C�t�nE��֝�+�E��|�+��}6
����s�U�؂8�f��-��oUD9�VD�yB�S3E�Q.�\�!��>b<�!���h�ޔ�@����^"���GHz���'HU��異���f&��~dӜ�����Ϋ]ZO���, f̡o&O�E P�:J	���@)1$`� L�R�c#�}�� hG �E�H����_��$_�t�3��v��g��<ժ�!�� �?:���b���`�w�2@�x>��g
�@��@��tj��$@*+P�UR�@���6��@��(
@�S��>�uX(�@�?%��>������'��|�W=�=���VAʐ��9ݵ�S������C/Y��r�����{1r<Y�{��E|>�ڭ���#��(��e�2\����WA��d>�!���"=Be$���S�6��au��Y�5[(�mAY�=F;��\>J@�_?[���J����F:��L��eJw��g̣�})��&"��E�).%|�;�/"���L�
*��T��,~X3�#[Q�����������b/����!ˆt���!��+���b���JQl�ȶq=n�gx3��!�\�� T��]"��.�ϝ
����� ��rj��U���o����=�~�G��m���p��N{Mr��rە������ '�I("�l�
c'�m��H� C?�9�^��^�F���a᧐ݥ,2Iz쓿! l�) ���*��S:l�Y�^����ؽ�:6l8�%r���0����s���Q ~fc �� ���
�� �����y��ݪ�����j�F��"�,��ǡL��rޖA����>������b�]s��s�{����z�����mHv��F�TI@����	�v�-��c�T�.E��C$�e���pf��	��;-�0�c׀h�zD�֫y�(�FE$� �v�S��er�D�mB�s3"][�ތ(�D{R���>�*OH	 I�#@P'z���12�"{��EC΢)gE�h�O�;@��1Ə�` �=`����HJ�G_(f��*	����INM���6�_�a��G@M	���`X��M`�2���%�)C��F�3<ȿ���oz�:���y>����(��F���4�Ҹʡ�rH�:�iU�4��l�@�P�%aOP҉Ґ%��(|��d��ߊB?]�1��]�m�����`��Q�P+�x��
r�;��P���c��3(��*�_�\V�9$۫�����U2�|�T��X�K>eB�e`�T����L��AogP2�7� U�,�	�	�Q�܎�6��פv0X:Q����Pٌ�`J�/?EE�%Mޑ��J^��|���_>߇�D��fy�� �G���l/�>$��т>ח!�S���<�:�5 ?��-Q�=U�:P�څ��'���AK� �1,�ۼ��_;C����^Ϫ[M�h����tr����>f(?�:�%��1��������	C�)�cYǞp]~,p�@I�8Ы~	bt�OU�����P���������C�0(�u�Vk�M�X��J9-I1��u	�Sk�� �K	���@��Ч�?/��{,��� '��$�:[�~����Q�_o�B] "q���Ǯ]W�^��p����~��0���۟� ��/��_�;u�>Պ��%��]l�v�!�5�(�����ve8�N�aݔCx�w��>� |�w��!�|��W\���t��)���R�_�F����&FO@����G
�qq�������Iugu�֩W��T~�����͠�0��G�u�)67jHդ�߬B	�U�l�bS�0[bW��۵��C�c��0���Rܚ�A	��yS|�Ԯ�H	�#('O�(W��Ff(�(�˩O�������L���f&4ˀ9��2���z	��7ˀY �Y���2���`�p���l��Z�@��T4iछS�ƥ�|�5�gOY�?���\?]�#dT�N����������`�(�zG��� �1��R����KK#�W�P�e��re��Lb#؇R6Xe����n�R�"�,�>DQh
)E��(�(�ns��G	�id@�#Ƿ��Z[5��&C-Ǉ�UE�f��R��ra ��0�+�U���A~@-rYm����>��R���h�y~��KP��`�;�!Kvp*�r[�� ˕a�Ǎ��!߷��^���VԦt��a_��H!��]�'h�f��>D%�"�Q�M?G��k!??q�k:�3����v�?���ތ~�YY&���y�/Sd��}n ��}^ +|�~AH#�oJGxJ�Ť4����'�b�_������~<�B�9�1�'\�4֜>f�=O�Q[5�y��+<������u�ןn��8����V��'�G( ������7@�5����5��7�_�Ӄ�R�K���7�1�%�Y���ln��Z�W����( �)܆M�!�e�]J1P@0#*�g[O	`qR�B%�픙B3��������򢞱��"U�.��`��H�1 �!�J �<
��
�[�`ݺX�`7fNY�o>X�O�:�n
����\ vL��{�~�w��.�|s�V5l��1V!N�X	춦`�G;����(�~L�X	��gas4	N����P�+��DZ��$�w��  �-A�C!/��>͍?�N�+�i�dW��;Y�?D�S+�6�=D�2��!�j(#U�^����R��˥�|�\+E�N��2�(CЭr�NB��lÿ��D�
��ёBp�.\V�&DQd���-�y	ޔ ߇H��D�E���ĕ���3E��֡��`H���f}3fD &��ހ������_79�����@�X 6�f`�?$!.a.��?���d`�0"Sޞ�0�K@�X�C�H/�>����$A2H���P�Ɠ�Z�>��$���e"l��"��<j���.EqX'e����}A����pkE�_��50��	E��B@�)���CP��!�� d���g�[Ȋ���@�`�R
9oL���P��=��H��˗�9�E�,7�MP�\���Α��B.o�y��(�ea��I|�ƌ.�d?�КӍ�<R�-���,2�܁ڸV%e�E��r�{�"ׅ������?G��(��+���Vqyj�\\��z�0�9�۹��
_U�z�E=@yC?������P����c��*f�_>ȪGT�.����Y�q�{"�芇\;F�׮���ާ�����	�^�K�x�a��<y�-"K)x:��O��I R D �("�F��z�k����/=T��J$U�8����^c�(����n�� ���P1�r
@�. �&�( �" 	&�@�1El?
Y��<'�( �C���V�5S�5����̔�HM �����G�ܺ���p��m��qE]`����������/���+S) ?�A����u���s��k����7x��`�gpui$n��í!��:�$�ښ,�x/E�����x����>��)˰n�I\?�ۇ��x<.g
�q��kr��H	��nE��v%).�q�*�M!?s���$;��Ir���v��&߬c�W��j9�/SH.���B1��#�|��\ �\�+E�ʿ�V��*�pz�b`E1��P��T!ء�NuJ�ڌh�@�����=ې��I>���ۅT.�c�>AE@�c-�Ȕ��:���� L<\pL,�� �^�Iv��� u��Q6vr�����ǆ��m ���� �� N�YKO ����	�~�*���!�0���(�(�痫��n .wEʐP�����E9��
6j������'(�x������S�(ڴ0�%�>�7 ��R���k��F�5���0��Y�|�ZV���)	��� +�B���%��JÚP���e�� ����k@0��*�>�u�������Ƌ�P���iE�{	��y�� �텽�(�C{q�JHq/�FKF'�R�Q�ͨ�GY`JY�{��������9�����g���R�ej����ތ��V�|qD�B�4꾢,�*b�����G*�k��Y�ј?���!��0ڪ�������ݦ�~�c`�)�C2�Dg��\?�Y�#�=��F��20�􌢿Gƛ����9�Z՘J���C�`�����-����X]�G_�}U����T��G�)n[�k[H�OY��6Y��m0s5#z���^�1*Iy�0AqC�D!%� ���vC)S��b�Y�q��У�r@`�9$+a�m��"H�����&D� зnyp����7Bq���öm��F�0o���W�-�'���^���� �����/����qbV(��������W��G����v��R\\��+�piy�����v���f��?~��_����3
�
����E���4XI��,���\(��e���~�1���H��@��#d�Q2>@'��	RܤKr�]�j_��Opz�8�v��?P�nӌP�FݨS�!|/U��B<���L�O���T|Nd��d|O���4�ϐs9�9����R>E� �W��� ~7
���VʀE�vB�T"�^z�y�����qmDE �������@��#��t"��12��$+�[��Z�����Cv4Üh  3�����ܸ��/���(G	pUp�0�m27�	���� %l$J��S�1J� ���`���q�ie6��P#��b#r�b9p����l������MJ�T>��)��IW���� �ﱁ�c�:�7�*x	pm��;�s^���a>4b����04zz�Z�xĊ��"U�4�Ra�K�Rr��S)H�l+(W��+��W��Y(��ށ^���)�yB!xL!�B	e�8�!�����o"SRr����@�]P�߬v��JX�?��Az
@� ��F`F�����d% 7�
پ媋]v(��Ŭ�	(��¿ȯR�UT3����:q?G�"�I/����b��+�vJ@k�S4eu�>��񭨋iBMd���PT���
V�(�B*��eb%WHQ(i�b����h��|,��,���)`Q��Չ]I�Q���sU�7�C��\:D�e�3p��>��=�o�� V��p�A����U"���z4\'G��1L�z9��iX�2�>>�K�y6��$cN��I
d�/�P���T��RI7���z���ja���}$�e����/տ\�:W��k�ʖ\_�пjn�r�����SFQ0(�s���R�@���>�9EɄ�P�$mʰ�n�u�}���Rr'�C��.&�M��J�VӌV������Ʋݍ��	@`5}J����	�y-�Ny����ؾ�2֬:�s�`Ɨ�w�?�VW�}�?�� � �;g�T���_��g����#|����͟b���0���X��N,!�__�/_����[���/��_���oWbٜc8�#g���ʁx�N���8�)��J@%�a��u�	1jl�*�)w;��J>��}����/$:?R��F�k��-���R��gK�z�.'��|<w�f��H܏�Y�8��c�:NNd��o����Lx����P.���2%�*��Z>|)�7�UlJH�-C�� 		p�A��Zĸ4PZ�v�mH���tJ@��d��	���K]�����^M. c��"0$�G	��ȕ��" �^(o�Ȑ ]����B:�"`P���UqU�H��Ԩ.��tu@% r�T2�1 "��Sv�	��x�//=�( UMc�����d%6��X�(����!K�� �Ͱ֓`H�4�ϟ��)�UYe�Ƥ!�n�zYY.�Nu�(+'J@�0�`�BE���n� +���n��S�P�c�(�E���)
ogX��8���(��8
X���:d�����P�*8����x�����H��E�y�b/`%^�𕊜��:�SS�/bE^̩ܮd_{��.��~�z 4`�W�q�Z��
� �K�pOv	�>AKZ;���!�"׌��TDԢ<�����VN)+��2V���T�3�ُo`ܮL�TU~u
?�	jS���I�V�_��o�d�?���!��0p}��z��_�a��:���+ׅq0�ǐ�:���p`��/` m�ꥸʺ++ �ZO��2HP������G���WPE���>J��O�a/H�4r�j,��+���ê�������8�_�,�9-�l�e"���� �5�`Ă9��' ���OzY�|?�D ��W�d ��ć�6
�}
@+���u:��.�p�� \�ٓ�8���6_���ٻ1�
��c���M ~��_P ���s���<;��� ��3S>����M�G���i
���,L���g}���[����o^��O(��̙�������8�+g����$�:��㙸s*.g�}�W�r�a7�i݄X�w�};��POT��1)�N2���2��>��Hw¬���V��}<�Í�q���Hq8��p�&Ñ���A!Q�|(	.���z$nG�5�s�d*�N��(���LJ@6���R(7��}� ��
Uo@��x��D�c5%@z�*p�Ю$ ً+�o�� ��( ��Ὂ�S@�ͷ� �13f	��;��3���i�����>iF�(H�0A $��ș�D��#u�L��HI�ʙ��(͔ u��q� "l�ig�� ��Sl,5	�}����K+Xid��I�ˆ����Q
F�`2`�MG����3 z��P F�٩�m��}.�zm��n(�rI/ Vu&56�U)�$Y�J�nW$Q��Q�ԋ26zel�J���P
Jb���}�A1(��PJ�:Y�?BI� ���=�:%�m(
����{�?���Et0@9���m^�W��"9>�����@z�Eih#_�	ea�
A@-���

@+�z6�M�]h͢ �P 
��tP���:V���R躪)P��h/���"y��fvQ�!����P߂��V��}T%��2�l������cE�	�]��A�*?�u��P������<�~=����o�z��u�׵6��)�c�u����YU���ǂ�+� W�!�325��	�z��I� _Wz���_��e7��5a��) ��2�;(�R��Y0%�U/?�\�WvA��r{�_.amL���\ֆ�a����տ�#�u�) �?�
��L�o��Z �����&�������$V�	]� �b֠�߫P�xܸ¢������.b���X��.L�|�~k1>}m6>���5���%���?b�X��&L{kf|2ӿ���_��goN�g��)����XVP.Z˹��b�Gk1��E��/3��_�b���X:�4vn��ޭ�8�3������$\c�Z���?��28����)�f`�[5 �� �e����c���p_M��*�n�0��� ��-ÿ�����p>�'V��G�`w0��,�{�a��e�'��D�h�������x8L���x�\��8��d
\O���E�B:�.e��jɆ��x�ȅ7E@z�ni�D4	(�%@z(�VJ�$����H/��+����b�0�C�(��"� 	��`�9��Q0$@���ב=�����P*�qc�i7|s�P.���H�\X�� W�C椻\�{� �)�'U�"��H@%�e �f�%��	0v�� ��=d�t2h�dPTVS�a�rX߸C�H��g[>�'�	P� |�ʅ�%�:��"%2�J���_.�"�'�QW�T�{d���j�i��&HDy� ʓP�ܯA)(UR�|LHq\7�E�)QOX�?F1��"B�@d�CMe|AYd'���p^����<)�}���\
Aq�}��A�GqhѪn"S�� �	�!�R֌J�C%���w#��L�z����ǣ�!V��]��t�{*v��j��j �}xPD��Q����!��A�5���G�����.JS'e�Sz�{U�3E5C}�g�h�Y�Z����4d��>�W���5�c�j�ns�!0n���� %`�0ʠ�uP*G��R0��D�.������Q�Ͽ��C ��WG�0�e���j��J�/N���&��)S���L�����5s��Rɶ$ק0�c�_�ʿ>_vQ1�s��\/)����:�E~�ݯo�1"E�EB0� �'=G�rY0��_���DV�	�HO�@j�$��SZ�0�J% nw�q�&�/��qW�c��/bղ�X0c'f|�_����a6>� ��/?����K��+�~_�7߾3�?��i�M���gb����s���c�˱��5�s�p\i��uc�7;0�͕������3m=/8�-��us(vn���8�;��'�ʡ�<�;�ө|��)bU]�J�\u�^�e��ǱnR]�R�2/���~A��Cn5(����pM��*�Z�g��r��U�f��@�O�����[�"a��f�+V��`�'�{#q{?e�`��.q9J	8�@��N�k�R R5��IȄ�,x^Ϧ Ho@�8	�zJu	�B�S=��m�ܳH���� �d>#�) ��~En� `�� 3�� �!<�r\�NI"7�$�H e@��JaJ��7P U�	`0J7��8G�=^W .�?����nL��%T� ���H�� ��E@���������.6�j��>6�"���������}��f�= " 2�����f��������.Y~N��z�L2 P�U-���Ъ.6���
�e�6��u�ߟ�A�@��^~�ŉ=(���S�(��SЭ(��bPB1)Pb���h
C���B��.EY,��FQ"I��Q�� :��ueQ�QIQ�� TpZ���b;P��ExJ� �Q � �Mx���1ow֎�Q�%`m|���4��1�U{���Bd����AO���S�J�3�-0���1�r��f�И7�d@¿!��I׿�" ��� ��?jb s�z�6�އ�����7� �����J��E��%��$U��>��_�-��n�駥�_�??�
MV���$�ep�ڧ�Y� ���G�
�j�?��~��2VŸֿ���`�, ������{�&vS ���1vL��:M <5�m��pꘋ�-/`Ւ#����& �Q >� |�/����7/�+~�����{_c�'�0���*��}6�>��o��S�2��Z���o@{[PZmw�3l����@9X��ߘ��36``�zl��͛���{$��]�t07���X�O�A�F�z��^B\D@B]�݌�g �/�8��h���T�;��g՟���?������h\�����pm[(nl���A��#7w�(����Qp8���p>�cqp>A	8�׳����D���+��J�Q����z�� C�� �ە�C���I���(	�s�v�=���H�AV0�>d���c8G��`~�\`��|�@.�`R�Q'�0�z��a�&Rt�2��� �" ��k�FGi���q�����BS1��l�(��"�g`���ut��Q�q���r�5W��s6�z�����]���G�*���7c<f��|�-'�����!�-�k�P���rz`�	ёeU2����Ʃ�H�1^B�O�A)H�E��|iʀBN6$��i���r"9�P��C!9�$�����x_)e���R`Av/�=Uc�c�2�u�P��2j>��7��v\���QՆJN�����k�L�~���d]����y���T�:���uJ��
^;���Ch-����H�'��Up70��rP�@cp�u�]
e�Y�)�/�ÿQ�/��Iz�Z+Gp�땜�G��l�z�:����>��R1��.���6�\��@@�O"&�=���ص'�����]1W�����K��A�����rT�s=SG�P8E�%��~���.�+*��֩U���P�	�����g�{��O���- 	�͈
�E��ƣ �Ni���ƕ�8y��w[c��X��0Lێ���o,����'��~1��& ��o~�[|���������LL��;L�l&�|>Sޚ�]�o���6�๶��P �c�#X��V�ys%�ys.�O߄��`�zo�u�}�qc �n�lő�8�[v	$���XI��Q� �ډ" =��JԹ|/W�`��7B^���/��/����q1����le"�'rp�h&��?��[{�p}W�RB.oǥ����)W6��@\�@��� X����0�>GJ��#1	p=�S�|�D~�xR </���j&�?��1�" ���,R�$к�P�P�*�;R�R\Z�ڊ8�H��@ �W���ϐ$Ї��~�1�) j�Ȕ�܎a���7B}��0�<���G�c�&
�A�����:EF6$��o���"J ���h`��"�\5(Z�"��T��E.=59l����]rxi�㔥��t�j9��q��q�Tu�@��v� ��lc�-W��IO�H����3*`��FX�_���}l�Y�a?�vh�q8�@�Y �}[(#9�Z�����ϯ;ʘ 6�f)	�E�H�t��T�J�@�\`����."G�������>��I����!b ��"r��h�@t7@��9�㟣��J��xV۬����ְ1d�*�)C�1��.Eu<����򱆴^4g�^����a���1���~D������u2��ly��v��m�f�1������X�+��\��+a�˺!�8&�2�Muq3�9m�c�A�ʝ! -�-D�����)���S3�-9G�}�~�v�6��,'����#c(��\��(r<�\lj��a>�uB�}��^!�Z�����>�}/����(��ud��H������H� ��Z�YT�O1��gk�gl���$���Bv9i���6c��D��(Y�U׿�ީu�ۡ���B��Bo���~p �N��ȴ�Ӣ�����A�=�{9ߣ	@
���1���$��hc D Q X`�ܷ@�o9 Ύ����	���ؿ�
[�Q j0������_L��� ��?��|:�0�����lf�@�	��וX��&l�h��S ���`��sX��n�{5����_��_pK6xc`�:_���zv�}[�p�A|rw����	�F�y(6��ǳ�p�2�
��t!�m	w���̻�-��<�=��Ɂ�)
�I�[�	���TXHƍ�|��|�Ѹ�5) 6�<?υ����镍�n�t�����;pk�&v(#�p�p8·c�~4� �3��<���������%~�r�����^ ���QD	(F E ���K �%���wk-'��sx�#A��ۅ$�'H&i�ϐ.��{�ڏ��A��Q��@�'�r] �J@C=��}N�T�f)�E�d�ȼ��e��I��9�M�pU�� �p#����ǐ�����&d׀qְ
6
j�t�K"��F��`Tel���4hRٰ���N<6|R��K3xe`�:K���8�v]�;U��*m|�XF\K���# 2@��	h�E�õ�@@] ���� |_6��3!�Y��፵�
�� Këz�������E�M0Ʊ������Am��H@�L������q��Gi����D��,�R�\���|��P�רa�\�׫Oau�S�<��{P��K�N-���4V�YVV���LY�v�w����%��W�"��DR��{>���R��'MDP��;Uǲ���H�t�K��a/���u��"P�ƥp�^ ��z$���i�|V����������a<c��N���6P���`��djF.O-���KNS���ȩ�Vi��}IO���w;?Ã:
 �_.��R��J�������+&�fA�9�Vߞپ�HuH.�J�'Y�*��;a�������8O�L�R�QLI5(J�������`�'��
���Ky��T�\J���$0~����.%��lW� >��" ���� \>�S��pP`�9�Zp���w�ŷ�/Ɨ�������O~9�?� |>s�� ��߽���ތ��' �f�����`�;k0��EX���u�X����y_�����n�.V���G���(��#"�K�58��#j���cٰg5�p2����T���?���wNdh�,�GSa}8V�ps_<��ŕ�~���-�8�1����4?˩5^8����y�E��F\��+[}qm�?n�
� �f_0l�����p8�� D��H4܏���T,<�&��|
�/ehp�@���	�]�`�*�R ���nM��	y�!λ	��H�{�$ 5���YA=�^�<�}^�0%��/�F���>M 	�`��7�?��U��.��PȀ�ȋ�$���Y�7�$qc�@Y2RN�X��oih*39e�[%��d����4L�I��Q���	�2V@�����T$@FK?ha5��)�jkZ��\�O�[�t2��8K7�s�U2��%� �j�@;L������W'ia�- G(`�ɡ���B]�X>+?�V�iˤ��L>@vp^���Zi�B�9t��|�*,O�w.g#�^��w/�E@$�,v��O� ��$JzzP'��o���P j%���JNhLa؋h�P�Ы��ԥ���e��5���0jgHuP�;yĀ�n�.
Z�
WJ �İ��cr�}9$O��'����\@��N�O�oF�q��(�f�x�d�C�J( ��Z)�)�a\@>��
%�����<�����-b�`������ 0���
�~�p���h��"@B'ok�?�������I����w��c\̧��� U���`�H�����M`H�AA�� �#�(H��<�\��Od���� H/ ���N$E��P�	�{��S`s�p��p�	v�����`��K�իs��o��翜���/>�
�~6& 3?���_-Čw�7Va�;[���}h�g�&�ރ=�.b����u���b,����Ƃ5�X����K�z?�"�(�6`�� ������qtg8N����}���\e�_;�*^NU�:�Mo����X"nL��|��x\�������k����[Cp��s������8��rt���t��U�8���6���zw\���[�qu�n���^J@ % ����`�(�G��~,�'c�uF�����Y/ 
�h]� �2E�C%B�� ԥ��H�v���R �|!޷�"Ѕd?���\�����!?�V��f�0ts�2�+�hP F�5�L~#��y��|���0� �%(	�c��vW�RPJ�PWS46U�O���#�Hx�{[k���
:���q�F��*ZvH`��&6����I(A�갑a�(�!�����:�M���L�r9߇���'����������}�!��d���$-��,mr8`;�6������1�u�#?��A��7#���V�T׭�8+	�"3��D����*�bc���Jo�ȖH��������a�����Ai� J��) }��KSx9Ű�ϩ�D%��*qՔ��d
��Բ�a�]�
�*q@!�k�q�H#?_�� ��Mz������t�K�ˈ�N�.��f��M��KիV�n
@�������!�����:�O܌�19����m�uH����>��~��~^9B�"�i~N,�z�2P�#�_���.y��Ea��y�ǩ�B�H�e9%"���o���O�4j��ADW�s=�%�� LD�'������Ov?��8�w��7�#��<^Hi-L$����"c�'K� e �: 'I�#+��T�ö4��U�=D5 ԧ�n�;, �G���:x��d����a��#X��N��h=���߾� _�v6���w?�1 ����ӯ1��i���LV�s��s0�KV��/Ŭ7Wc�[��}Z����w�%
�^,|w-�����m��9�0{�]�[�EJ<�`����������qc �2�wlƾm!���pdge �2�S�g ��w�`_�N<.2��3���������魁8�9 �7���_]�<qd��r¡�� �X���qv��o� x��6/\�鍛�}4	� ���'�C�r8�����:� �s�$�������@��( �Z�p���U� ��6 ̽	�h�6��t ��%��$��1R(�\��^��0V�c~?W`gG� h�z�w ������o �>>'��͏2Q�m���
�>�|��E2P;Fi��Ay<�h*J�Ill��C�d6A�IZ�%�Nt!�×T7y�VQZ�FO� �zVqj��TLl<�)uִ&���bu�.�*Yy�~|�����.c*�Or���d�Ni� C �9؀��k�3�T��j��F` U�c�.�~_%���ve��lJ�׌��h�
("	���w�FW�n�������P��Q �Ỳ/(�%Q"C(���A�Q�b�{𷫈�{�Q������j�F5��f���]���(aHM�v5����4�7k���Bik�ot��&��}�pmg�v��?�.�MC=���pm�������m��<����a	=Y�>42͘��g2��4p���(�,��^-|O9J@C��?�O�T������ �70й���\�4���a����(9$�uԕ���F�/��K��]!��_��Lm�0&���0S��L��)G�L��11�������� ]&
@a2�:I��K�EnR/r�AI=�>W�Ȋ�Fz��D>BR��5"ܷ~n�p����1�v6����vl_u��R �ى9mČ�W`�ᛗ���_���' �) ��ۦ@� �P �b������V�c�*W�]끹����Ῐ,��bU�v�?6l
�6�ss �P�oŁma8D�n�l�4!��p�duop�w|K��5�mb�od�o����^8D�8��W���*XiOn��
;[}'�:��Z�[��qi�;�nw�x*	���6��;��@	p>
���<�S��:�ﳩ�>��KY�2� x����.�?+�@#��k�R�`
@( ܳQ>m���@���h���2��0V��H�<K��%@�		0�	~K c
$�t�)�k|M�@��,��lL�S��*���2�!�겜�K����}�j��tk������2�0d�'��4|lkJ�����,�ꎍg3�fV�έl��z�2��
�.�U��5vߣ�r:`V�|��@z D ���^M����H	�Z6�5�jJ�x�
.������b#^����f,����JN�Q�J~'�V��7���e	CY����� N�};��3%\w�#8���o+TP���^"l�{�*�[5_��Pũ����m�8��{���sȘ���u8^��V�����f�߫Bk��5|"k�{* �z J���o˿W��Q��JWO��߉�:�����(:r5�z>�@�j�w�$=��2�P���zd���4d�!r�]�PB��\����^*�qȮ�I0�ٲ�O��'�.= � )����7 .����\�C�N1�?! E���~E�	�]�,�(�l#�� ('��"+�Յ�v�6#§���p�����bq�L0�p��m�ع���=�������6�x�kK1�w1�_���7/���E����X��vl�l?���= ��] ����+���q�Xt3��`������s��b+�������9]��׳B��J}+�`;e`��@�����_��zN�����:��2=�֛0�u�u�>��U�ػ�{W��~�-��ƑU68����:��zg\�䂋�]py�+�����]^� oX����^��� ���H8<�E��D�N'��t
��Q .fjpU ?
�/�G� �*��M	X�:T"�n�
���
@�o'�d, �_H�Sw#;�vĀF^�(
$����' �h=�з�-��0�sI��|V}:/ �P 
�cf(!�"���!2M$T*��(K�}Ք �@���JV��/`���2hظTm � '6a���:U��kUಁg����G���7+�Q����ۥ+V��>`��.��5"��!90x�>��Vg�˳��o! y�f9Y+�&y_�����!��g65
6�7��a�UK�q���.^i�e �P��"K�*N;���ߛ�`@�jY+��w.�/�>���_�����r�]9��VH��d*����9A�^�Z�g-w��~�Ƽa�j������2�]!�.Q��e�I�w���)��]�0�$��uJ�44w��S�uD��1�q�>��ep�r��z~o�����y\��(B��H��yD���q��KB�Iw}+���o?��:���K��o�|�Ъ����~�JF0��8N ��L�ɐkt�1$@��i`H��� ���� y�"�y#�Kx�A�<'I�$��S�ų��{�i/���QlG�:ЂH�:����v&�P n�ƹ�n8���V^�z
��o�`�G[0筵������Ř���?7x����`:�|6�?��?��y_.Ǵ�( ���w�bۧ�p/����m��?��p K�^�Yo-�������Ø=�3��w��1{����|�+��(��HX��k}����l�}���cٺʏ�b�J_l_�+�hf��;�z;Wyw�^톽�]�W�`�*'�Z-8(v��߻ڎ�`��*+Zc��kmpl�Nn����qa�]\�挫;\qc�;�v{�v�7n���>?�=WJ����GzN'��l�) ���p9W�p�׋p��J`[� {m��[B<�)4!ī�^���mC��CD�w�.ĐX�.��H�}��g�
�Gn��0t��Z�t.�w� PTO��ɋЂ��Zȿ >�H�O���'����1��g@��I��a����b�X)d�#B�θ'B��K1�Cl�����6�d���4��nW�e����9ِ�T�Z��b|�f�^t9�Q�S���[-�	 �GG}FA��R٪� p/@���x��EX�Bi��PB9�B�	�<�]Il�%�)_�;��h`�C���@~��~����{���K#?c?k?{���˫���#���6�7�-�Zn�����r�X�{�4�;��g��z$�(��e^C.�+�k�&4��ԀB]�\&u�"��$��P=�M�NN�<�\��z@d�6�����WW�a�l�Tn���jH��ɐ�t�)�2��-�zTN�,�`kp;�w$Ⱦ�II�9M�AY
���v	a>N�7(N�P�4H���N�,��'%P�*�ql/c{��ia��x�>t.��]����@\��c[l�g�el�s
��a�}���ڈ�Z���_��^^�s�W��1�� -�|潿߽��?ل���CGf04� ,� ̘z�;���m1}��[�Y+�0g�;�������~��K��b��X�U+��f�7�.�ƺe^��z`�R7l\�MK]�36-s��e��.���w��+�b�J'�H�c�=�����߳�?�*k�]iM	���5V8��Fq�pz�=�mq�EJ�eJ�����6��`���{}�? .��v8ǣ�u2�g��{N������� V�A7
I	�n�!кA��C���Z�j���߄P�O+B}�!��"�;��P #:�1��#�$�ic�����O��2<Nr�/ �0	y�;C �U�/��
��ɂ�@s����	)�C0F�t93�d���
��j ��
Vy�CD�!������ny�V�]�̚��b�.���.���x9ِ���M��s[�7��&�N#_s20��	�5�?���.:"��Ҡ˥���\��p?U ̘�
��C"J�^�a���*�"��Uw;+Z.G#����n��uV;Y^Uղ��Sٲ2� 6��Ƃ��?�/:f10�?C:���{��#=�yՙ-)w��>h��{\��`�J�b�0Ҧ\G&C���@��Xod,�ꭐs��(������K�T����O@v��uR�|Q�@��. r�1�8��N�~[.+\#�����!�H���X�F;���&N��au"��y���;ؿ���9������wc��[��/0ﵵ�����9`��s���EX��|��b,[w
˦�E{J�@z �~�ӿ��)s�0u�%@v8c�JWJ����?�[㇅�E����_�����Ɋ��X�ĕ�`�g�Y|�8a�bG�Y�@�v��_t��Ɩeز�[V�!��u��1����w������M����V8����Z[�9����	W��X������}�p�{<�EP bX�'��B/g"�Z6�?�7|��V%f���䰿0g��G#"|Z�ۊp�����D>DdP'����1$6�	��p�}���*'�}��@���\�Æ�>�|V�/ A�>��c��d�@^o2
H���_�����_�\G�&Й:�r�!���!��|�B99���D��_�XPF8���]B� 6��ҍ�Ƹ����G��V�XH�.h�E ���+�������I_C�3�(R�7�Vq���ԑ�	3jW���C�]j� �G����ˮN.�P�l2�'
�D���  "f`��	��JX����|�\u��V��P�,������\9]�vFE���bE�����	5v�������$f1��㯃?������\ߌ]�#뜌G�ny˹
JY�(�� 9�As�%�_�� h� �����VS�-�j�?�d�}�&	��R��X�=��>��ol]2#��.�CW��C(����X��$j�����Z5��E��d?A�o;�=X|9V��*.�aw<�X�����oa������I��� V���^ߎ%ڊ�����YS�bǆ�� ;w��4��ϗ���P,�n?i� �{q`�u
�A% ߽�gl÷_����( 7�����ӗ:b�
g�\��V{b%`6�%`�jo��`�
,X��-ܰx�3/r$XJ�-���w�l�mNoc%Y�ЖR`�Koc�[l\f�M+l�y����6�����/�g�-�[{�Y+8��'7�Vpn���+[�^�����]^p�㋻��z8�G��}*�g�( ���Ɋ?����P�"������z��*�k�ր�fD0�#�#*��a�t:I"C�'|�)b�	 N	���LH��FZ@҃z�ҏ�099��
@C}2r��tr#E4�"D*Ɛ�ԑ���(fPct&���3 ��'��A1CH�g�~m�DCZ�,c���r8��P�ٟ�@�}窻��iTg�ҍD�"��P�x~9����S��g��̠oQ"��85P�?���oND�=�# ��X�����e��yp����]&��� ux�� M�d��,�� ���6	�����%?{����g� ��L.���e?���oF}����ꁯ��am��=�s���g��@��?��Oj%b©�I$�� =�v�ډ����`�
 � ��|r{��"0y�:���g��ߧ��	KRE٪�����$�_�ￜ�6� p��` O�d�O�( �◁��=b�ߩ�m2?'��RI�:W)����V���d�W����핂�r_�KIq(% �2�!����k�Z=/d��X,n�ąn8��f�����a��Ǳ���X��^���n��Ӯ�� �[��Wm��/fc�ؾ���p!f|�s�܂�_�Gsʃ�������v�9|3�*�YpSYS�1u�%�3V�c&���>���3) 3Wy���M���P �.v�<V��:�;X@2�.����vX���B`���j�%�k�Xa�2+lXa��+���a�����m�5�����+oa�س榒�Ck��X���p�pv�=�or���N�J	������NO����c��(���C��d_�b�g#Ħ �wJ�PN*�X��5�`�G1���Q�ҁ��G��z��Џ|���nDFt#*��ϡ Q ��tS z��ߋ��>J� �vY����ʞ�B&���1dw�A�^����k`��I J��3|��(fc��Iw6tc��
;i��P��TìD� 6��w�[Y�Lչ�Ґj��tӲ&���1.J����2Џ2`�u��(s�& �o���/��aQ���@nk�k�|�~�j~�*6���! /�P�[ ��`�n��B�WUzr�bA$��M��C`�T��:US�=>ׄv�Z6�"{�[��<Pp}�����G��5ơ�����&J d#���pJ�n A^[���C�HԺ�zD
��J���p=7� ��] ?N �Q�14)���P���8�G�V%�7ש�����������i-׷Bۈj�5lO��y;��C�6�ە�V���!�"��1�]�{���v�����Hlv���z/�^℣�m���k���yl{���u[�8�M���
���g�ʙ�8��8�/�cє5���_��8��Ax��v�P L߂��؂���3/᫹�(7��";|��S��Ŵ��N	�A	���Ӆ�^��^��En��ș8`��Y���l1g��̳��y6X8��Xc�|+,_h���m�f�-�[z�ߢܢܤ��e�����7�Uױg�\sG�X��:[� ��S6��.�D���f������~?
@  D	�߅x^NA��,�X�"�v!����\E��R�(��Wb��#6������D|���=�yNz�Cx���g��?E,�^ �Ѝ�������~d�"����\
�\ ����9����C�l&� M��P'�a�#c�q�!�$6lrYT5�[UjV�Rk`C�(ݵ�z6�ul���*ԫ��0�^�S_;�¿�����@ d����=&�#��}J��5l�� Pd�-�� K7�$ �]�2`��!]�ɬ�(�0Vi˼ b0��3T��H�����R�K���^{�l�:��c~���M���@�&���d@�1"c��Đ�l,���yf0�@$@����ơ�=D�� ��O�d�/ș?��_���wXK�n�܎-���T�����{-�	�Z�u�ZM�֦5�]-p�"��o� 
��!ۭ�����Q���l���;V��p�Ytv�3�O���o���W���K����}���M ~K�0��0k�lY���{�r�*�z	���t{><����`��_}s_θ�/f������6�v�m|��S�;b�rg�\�ƪ�]�b��/��n������.f,rČw0��9��|G�ε�XQ��h�-,%�Ya�b+�]j�u˭�~�`���� ���+�cٱ�vQ ����z�I/ 9�����������W�:��������=�p<��#�8
��Q𿘀�k���F�]"��R��*D�� ֳ��M�����|�C$Dt!!�)b�!!�9�A|B/��׋(���nDE<AX8	{��PJB ���=�$��;& �C�FV���ȦL$���6��)o˼�Ms�(JHQ�7�pZ�V��������ۤ��K"ٰD�Q*S�~���I ���Q�@b��j�4C�,iH��iPe@PզTkDFs�ʾ[6zr8�\2U����Ⱦ[Vl�}�lT�W��4��K�l���1��0�}�����܉��	�ߐZ}����Ǥ����h�e�4�j l�j&Xl`�{R'cb�Z���!������F[n3���dArҠ8�g�$ f�]Z��ظ+T�K��Ϡ0�A��7�7��S��f�T�}���rX��j�(7rxiy�H�-^�*d�T(�>W{>JHШ�r��S�}&����I�;�@�^ٵ!�D.-��r�!ut 9��|��q��h0�� c�����٥���Ҫ�!�LTS"��Pg���0��:�O��� Z�\�
����}üL�J�6��:Hx��Z)�35Su9a�%'S~G�]U9�d=i��ޔ4̌�0�n�X5�7o�����)i����ߪ��c��F��l��nՇ�`.s�09m
��(����U��3y��������ٌ��U�?Q �}ip��5a�Z������TO\���p�������N?G����_���C�p|�	̛��ĔW`�;{�e�6~v��/�X8����F|��q|1�>��,��sS���0����eN�A	�!��f� ,��" �)�) ��9߆`C��<�����XD	X<_$�
+��J���VX�\v0�Y�Z��Pl[y�( ����rx�-[g��k�q�pn�-.�����Mθ��6�\��.�}�~�>'C�.A��v=Ѷو�/@�s)��*�Q�x�z$�4#��� )!H�`����xV�I}HJP$$R)���~���g�F�?:��Ѓ8����x�'p�ԇ��EZ� 2Y���M���K@�_�ƼbB�� R,P.,���{0��6����!Z�X���&���e��>��_ЮL��_;ݰ6�l����rc�����V�D%Z�ƆSzT�i�������1�>}	�	H�װ����ɩU�SV��M������`�1 �l����d. 9+��V�`� c`���T"�VT��ʎ��P�Ч��h� Ԑ�8���0��0nK�kSM�_9k'|R� /��e���2��0�uj���P��_>�������	Q������$u�	��(�n�.
~���\��ɀFu�a�&rt��'�2��$�*���қ$�Z������(�s�r�r�)9��P���7��
q��-��*p=�.�O2��S%�C_�Ч*�I9��,�ߍN����D��3�-�$�%��R J( %�n[%���@?no��/��*~~W���4�Vn��(���;ߧ <���F�kg�w��2}(p}�����m��EA;ۭ6�}V���8����-����+�՟ߗ7�Qn�w��n� �F'R/<@��z��+���x�M����/�ݜ@ܞ ۙ~�����?_���L�9z'��²y0w�z|��*�x� v�����o��`���|���c�|�Y|>�,��sS���t�����ŷ1m�#�P �]錩����J��O� L[��K������H��v����(���b��S
�P �-��U�nb͒�X���-���~�;�lZy[d7 �皛س�&�������膛8��N�����pa�m\YCX�[�a��wwz�}�/<����t0�.F"�j"�R{'�wK�^��:#�Z��nCj�C�Ev!=�i�ϑ߇��~$��a$qI q\飹�� ,��a��^đ��^D3��+��#��$R��z!H	B:�=�!�Cd�\V���GT/�$��:Q�|�߃��Ԯ��:$��_h&��A(d�El �j�;��z�b6&��wlD�`@�q)c$�%�% K6�el�����S�� �|6f:UҀZ`��F�{]��l�ǐۄ~%{�j�A��߳�7��fC��g��U��*�n5��P�������eW����A[\ߌì$D��P7����^�� �FTGZ$�L�!4!���3$dԶ
r	uA��r�ڕ
5J�}��Z(�����P��d~�I�e��a���E3����(�畋X��J-�Yo�u�RHu}~�rĉ��AF�+Ad��{d���v9k��:Q�)�S �y�A��~[W�j�S�6m��02���-%�\���Be	���/��
�#e�|.#�iY.�5�˖��%k�BI�Fq��t~�i}ԩzSe�߆"PH0(�ȡ~U���)uM�6s����>i#���u���E�9�=�N{I�W5�}}�n{)���{(���F<��I	$��?����G���k{�=<(.#h�3���=(�؍��]�<؆�����T���\U��e��_��E9𛟅�yY?c�z&�.]�5��b��X0u%f~���܀e���Oϡ&�U	�3�0�u���o���7�R 6��7j0�,>�q_;�o�����1e�����oW8�U�>�_� @�+!p����3��I���w�-�qw0��s)�(��J�6�
��Zc�r+�]a�u+����������c�5v����o�5m��rl�-Nl����v���6�m�Ǎ������=np;L	8�����������@�c>"]���O�oFb�=�$�v )�!�#i�1O���q=HK�GZ� �i�Ii#Hd��:�XR-8�rP� B��އА�	%���DI��P
�"6�	Aϐ܃��^���#5b i����I��Y�CȞ�\�.g԰��<_=�)�}��W�*�J^�����F'��e>Dq�Z��N~߇��q�( ��R�j��"`����9=��&���M	�6沟��r6��8HŤ��g��BV�l���VI�%��
	i6�U:"R�[����Q5�
� �d�_�ׯ,fC��U\�4�dVo22�$��F�,Ib���-��X�Ї��^H�F3����3����A��a4�Ϳ��P���	L���[������%��'�Z(��P�l��1
IA��s��( �ܮ�rP
En&��rbP$��2'�m9�LI��eI�})\vR,�jW*`�&�J;��@6o�:�b(Gh���x-��k�L�t����J,�.`��$� 	��V�/��R~> ��\?���y\"��\���2gsy3�$��O
���r��g���\�'��RJ? ��A�˅�(RM��c���=�:��6���_/��~w�٣�:�� �p�%2��0%v(����(�5�)�}l��f����c�϶g����a������� 8��ٮ�7���"Pz�1
�v!o�Sd��BƎ���ց̭���Ҧ��
��ϧb���0㋙���,�b�;__��o�O��&��" �f]�� |�Ŧ�	�W�/Ya��_h����`�3�-v��E��Xg�Bw��pw���w�l���sQ��w+�:b�\{��c��s�`����8�6Q6/��-K챕ұm�=v.���ew�o�=�r��Վ8���68��Fg�f�/�>Ǫ��:'\[瀛�`��w�:�u�'�1���#�+�+i����8�$ٗ!ŭ�>���oCvP�C!7�	��1r"#7�)�n,�^���OD�\��9$�P:�DVO�lT�cz�����p�/�f����׵~�ߥ�rmD�[3�ݛ�тH�{��h���MN���$x�#ь�F�w��(4f�u&�g��I��'�>B�_���,WIT<��n���9Ѕ���c9�������1�##��$��3dFu#+��1��>Ef�cEɎ���Ή�����'=����y)O�(>EA*Ic�!�v#�ӼtNIa�L�$�<�/�ѦE��(��(漠ns������{g���9���K�K���?Bf�~��HV;��{��ЇH�@��
bD� Ϳ�:2o�*��/ -��)
mH��f��{҂Z-��LJ�+R��O
�O�6b`,�"���2���Є��r����wd�2�1~����.dGw!'�����I$�	��{�dt���S9��\�G�����9�
�S ���L�v�v�3���NIY_S�ߗ�=cOd��/�y��'(�⺕����u#��HjrS�YIv2?{�!�$3�!�o������"�߅A$����$5�����>�o��)�߉���2�E���z���gh����r?�</~�ޒ��+#�=��Ao�������>�U�JRч޲^������~�����۽�}�����~<�Dw� �f�i�0SN�=~B�{Bq|ۇ�l��Dkt������_�ǜ/�b�{s1���X��nl��(*��z�ML�g�]���y��jr��4 �R�]������[z���q~��4#�\"�7 �|�ϙ����{�q�j�	���t��Wj�v��W��|�i��u�9$�Z#�6��j=
�բ�j-�����5��j@�]3�o������:��҉V�'����FmO��j���x[�s<��=V���q/���x�G�푽h��mr?r �H+��ưAd�>EX�cxG=�ٛ�ر��(-���Q�X#g:����`�{�]yG�o�=��vP\㈃k�p���P�O�!��d^{W]Y��j�:��7S��tk9��G��s#��c��|>�]���G6�o,x��F3|�&����=p|���'��m~�'��ۦq�`��6WN��|�v3��S;�pj�xN��4N���pb�+N����}�m��^w�=:��{���'��c�\pl��������o�}[���\&޿ѕ���P|�n���c��J�u��.5�r��zm*��9L9>��������#�~�&��:G6ܱpx��I9�������v����=\���/�,��QYn�O>�{��n�Ϭ�����i�ؖ�8���V��悓�g������ӻ�pf��8�Og���9���h���Ȕ�=CN��\?N˺����3�ܵ�\g{��v;㄰��u'?3?�1rt;�i;�M�;Xqzl;�:sd+����~�h�,߁Ʊ͎8���	'���q�)���wx��������t
���QQF��������t�����}�C��a"�Ab��Q�y�}�����5��!��O��k��k
|�y?K��/���S,0�����Vb���1��5X�����8�b��p��_�eX8m3`����6`�Y}�fϱ��=IȻ���Qmӧ��@�� �B�� ���l�� *�zy�Uv��洖����f�����ݨnu�.�~�Z�~�Z�ޚ���gh���wƊg��>�s��<tF��0���Ð������r�i��݆1�5���p�"�\q"t"y;Jc$��l�)���L��e~D�c��Ə"�U�oT'N_M���ع�
����XL^��7�u�l[p��7����Xx��®ŷ�s��I��v��,!��;x[��]��5�>���LxLG��ǌ���m��na��,�Yl��vص�ϟ�n��.���u^��evػ�,�M(TK9/�-��>޿o9������N{�a�طR����_eGI�k�ѐ���|��^a-�f� ��֠�)�m;�Yk�=k�4V�s�����ܽ����"V\���Ԛ��-�d	�~���[�ή�k�c���Ku&���:�!��1�R�_�An��?�<煘��=\��=|�=������N�^�u�3�nb�2~?:��u�;}�o���ވb�-bK��o����Z\G����������N��y4���5����q����\g�s����b׉}k�Y��3�۷,�]�eZy��;$2�+��
Y�	p��,�Q��:K��\��/�����J;_�ӫ\qck ��f�$����c�0:LFG��l_�����m�?��`X0?�ϗ��?�q���QGت*�<"������tP!�9B[%2/a���."����}�7��_������[L�l*�>C�p�K0��E�UX��6l���"k�}=Ћ��]����R �R �c�ԭ�����t�I|6�<��A�\�l�g,�ŵ��(�{�J������(E ��S�f�A>� �v՝Tߖ�è#�6���㵶��OD�2`=DAq��m��Ɗ�ps�|�>��6�� ��2@�+m
��0�;w��q�A?���xȠxw���}x��=n\񜹾�3�=����jc4���dQ\���`�[��r��X��" ��'�2� 2�>��8y-^��h;��Ml�6���Đ�ߺ@c�<J����7;0�� �4�}"Ҷ��H��8v� {�P &AI����`���OC�Z��>��OE�xi���g`�\��d� X����]�:濷 1�?�
�d�Y� ԙx��e�������w��gppC\��� �� C}2�$�Zǿӑ����S�kp�a?�WSHt�:(f���2���Ev/��L�l��{�\�L�8 G(�Ǘ�ũen���7��mOR�Pٍ�:����,,E8a(�rcDG�#Z�*����i@.<����X��l�h?J�j4��ϼ�����·�`��˰���W���T
������0��������\i7B�#2Ї��9?G��3Ըv�����0�)
U�@��j��N�hbX7:��i5֣����u���c4���ѹ�n��t����k?Z�z�lߏV�a2��з�΃hsg��ۃ6�}'��	%��[/:|��o ����{Y��a��<�i,�q$�+����!�'���U�1L	h��CB�S�D�+�N\�S������ C�`� ��)(iX���{X�W&��əLX~<�I�0�L�)L'���,{W򾟈9�w��̟K�&v���[�'ٹ�c��I"?  /bb��H��r�
/����5�a��\���!A��B`�oz3ߌ9�w-�na����*L��h����P�-�M	�ǉ�wqn�'��
���8nJA�2�:��%�z�Yo�H7;�_Jm�J�������B �6���������7�ooº���$��2&� z�{�9�zO.��
��\���4�X`�E|��E|�������vU� T�����
�0�A�����g�-�H���{ߣ{v���0��k ���D �@�]�`A���Q�ݓ@��;�����9��U]U]�I����=�Tե6|�������%jW����g��]+�i��3��p��Z�m�U̐_�MG�P�������p��s�;��o���Y���8D����h�x\ц�;��vx��/״���6<�؀f������F������>��V���F8m9N�e���^L{�� �'����/$��0��`�W<ÞCM�̟a������K�����Η�/� NUhC!P`�+M%1 !���/@�t �B-E�I�z�	��N
�@-�0��r���鲝�R��a����.G��;���>Tt�.A/��H`�����??�>�u��D8R��9��u���M�\���Ÿ	�t���T��h_n���N��:��.T+ Ѣ�_�r��U��9�o�D��+��^�"���A%r	��wCH��HpZ�t�M��؆��G���{���ǡ���\�Ͽ{���|!-��Wt�+z�  ����.`��1 B tg�A����h�	̴�a0�&�`3��3�qqOU� �'�uJ0�&�Bo�������B Lӡm�-�� q�\
�ե�x�8�/���z)+w����-���ne _[�
�+>0��qm�;4\`���-j�Q�c��~�^�j�+�-�k����<��dm����﹮	ז�1 ����5^a��j�ΊF<XN1XAX���<��,�]����67���p��픎&4l{�u����Ѱ��?��`>a����N� `��ο=\�x����QA�(���G�8�(��E�hھB ���GDO@ C��&��XE 	��2 ��Q�b?�P�_:eD]��R�I�
� �ôK�w��0a�"���Y(�?�ϗ#�����%O! �8B��"5���TwBI�}�" š�"�E��@Q�׼.D��#�]y��KA4�.���"��:�~)��O����g����_E��(B]����q��Ǟ�d�E8��P��!�y=2�6��c+�x��j�3�tۣ*q*�&�m}�w�����|��vS��kkdC)����� S-K�N2��8;XN�����]�?�I=��q���;Ag�,��E�a��) �R������$ ���� ,kC��7h� Ԯ~�16`9PU�O�����Yގzq1�u�ZٌjV�Ք���%-�Y�m�2�K��v�{.��|�ō���xu�w�����v�]Ո{����pg#�.���&4ߊ���J��z4�Ђƭ�v�M�ޢe�;�0 v�Jw�*��'Dy�'�ar���US@l{��Z��8��(9�	�G���ć��߁7��>��	T"��pw$�:�C>��jPI�Ǆ�*����F ��N$d�*��ȷ�0��U�3`>e����r7�ӣ ����$��ˑ� 
f�ڝP)�>�¥x��Ȼ�E��B r��G`p{�#�[A��}"�)
j��U���w�α=��w�ev���PI�����|�%X��W#Ź����Q�+}O�<�,v�]š�u�)��i��˔��lE�7����� �uQ+ &� �h[@{�)����l����ܮ+
x\�X�N���8{h��� �v�,�4�1K��lVG
8�E �Ā>i`+~R��!���|�'�_���x��O�ÇKM���%��hB}e�|�������F<�݌;kޡj�T��G��V��׀'x��wV����z��s���U� �5�ޚFI �li����Ā���)�9=/�^^�~�����h�݂��4^jD�f��mC�Qr@�'�g@u�_%P�1��p;N2�wnBŉVl� l� l� �� <�%�xQ ���S	�$l8U���t�ǿA �2	a���t���T ��W�����:����P�}U�e��(�?�ϗ�OP/ by��xo����� ��kثP�����9�V|n:��̕$�?7?��K��+��I���Z��m(�މU������\���8{5E��lO=�]jF��vE '�b�����U��-�����@��`J�@h̜]M=�i�`�95�a�i��F�i�����﷝G��v�y�����]a8�
�c`��
M�@L�_��F�4���\̢ �/CZ�	\*mdU.F�K���(� �q ��P�
���v�����M���F<����Xɋ
�{������ӽ��tg�3��z�kŊ�n�je���١x�=]��m�KT/y���������K)���	wV�ǃu-h9ߎ'[����wh:׎����MEZv�=T4��1.?ۄ7�0�\o�6���cZ~hA����H�� ?!j�M������}�h9D�W�:����{����-�u��Ў�'Z��x=�3��ӵ~lpT��̋x����.�l}�x�
��/�_`%d �c�`� PA� ��KP�����W�AP�� �I`��s��B��e�Ȁ,L�!�Kz �|G��璞'ȟ#G���ҵAW�_�� ����f�M���T��W>q��*	�v��/!������X8�[%� �lt�^�� <e��z� P�%ѹ��}0�)s�;�pc +������Pw���I�&��|"�%9T��*���^�(��vE��wC���b<��8�IҘ�rd{lB��6����ʀ��xA��Y��q�Q��
O7������ڀ�6��7���������8���-��M<��J�������� ��s����9�Лm���0�c�q:�9\z�`4�םB��v<�}ۙ^0m�Qf�3Z���9��������c����Y� �/Ej�q\,iDuq3%���V�i-E��_��-�lGͦ�x|�[P��*��A��f\_тFq	�5��\֌Z~���6�*j��RJ�/N!�]*�x�G[�rw#�-}����ۈ+����w������֋mxPQOqx�g��Mx���W�2�Ԍ7GX��ԄƝ��������l@;�}{3����g�@%b���uoqp��9ފ�G[��B��D6�l�(�˵��@�Apg {��TI�����"�{� ��� u�/���1�f�� ��U]�	� �. ����9r��+l�e�����ԅ�@ݶ��PC�_���w̦ ����@ �F�>���퉼��	��sI$�Ѷ�
PJ�4 Щ��K���H	HuY�J@��f�ymC��.��>�u~��9�G���}a�8wU9��xs=����/؆�����vŹ�R�B
��,�8�k��u	� 1��S�@w�	1����4��� 3�����0c�.�ƚ�h��gy�j�'�F�@{$%a��ρ��f��a���0L�l�ThXfc�}!��J�|�Kޡ��t��v]q��5%}
@ͪ4�[��fx/k��Mx�c+no|����Z��ZQS�WV���FԮ|���UR�ۅ�(bП8���)�v��yEj
^���Wh:݊�^�F�3�^��ݩ�.���z����P�*� z���[� ��jǻC�xw����t�&z�bd���s� �z	
��n���-8���j¶#M�����O���T6�h���c�v�� �� /"$���� AǼ�lIDO���( ��P��`$#��H'��@�<\��,_�}]O�\. �(���+��6]a��ϋ
u�u�����t����.�)���) ��!�D>P�� �'��>><Љ|�� s) ���3����WW���|� yt"���$ �>����� B�l����PI�@�	X���(�+�L	Hw[�L����@��6,�ڃUއ���46�����*	���#��z�k�/{�wgX�=kG[3_����oW\�G�9 � �� �H?
@_��;&ڎПn��Й͊_S���0m�tL:�G�`�pS������pӌ�������50y�t���a��&���t�h%c�E���A׮�A�S�\-i$M�S�ZP]܂*��&�2�OP ������K��.��Ɠ픂��.c@_mƻ��Q�ӟ�i��x}�=n�l�u���nq
 C���t��YQ�[��Z`M�S<��-���Z���\{�c�Y+�x����G��|m;ެ�}�oB��v��ư��~k�᪣sֵ���T��?ֳ �B_z,�1�m��Y����8�����a/�}G�) ��q� l>^���) Et*�������l(�����H�D�)�8e���(B=�P��`
��� ��Q��u�/��( ]��˂V�ݑo'G��.a�|�:�ϑJԽ�B D�*Pwj�a��������Q�%�q@���l��Ah7��%	��'Cu:�<XU��%ĝG�|��p����o�Gg�wG����~9aNx%���T�O������#����! u�:  �i	�)��WPV!ɹ�.��Z�,��V�"��X�~ �<OR~�f�s��W����p6�������S�1F�C;��ن�m����"��Z�~]п��@X�d�Lae/I�!fL�¨�0i�,h5��V�DW��6,�_�a֘2L�M���S`�K!�t�D�hL�O�,��0O�T��&����ӒW�\�@>��PU�@�W/mFͲ&V攂RqI�6��@U��"��s;��5��=�o�kc�ގjAu)��T�+o½��x���f��.}�ڼפ��P[t���ps��^��J�qk�3�7�nY������v�^����m�h�Ba�܆�{�v�	-G>��Xڎ����=_H�� �~���p;��W��±=����w�Y��;ъ=��wQ���lA ���\��� � �x�w.� ���u�L��W=�M ���t��>|?M� g���@Tx
�u��L�C>XT��~�{TH�?R D�3�?:P�%h�U�\w>�P d�+b��Ȼ�����|�~�kȻ�� {_]��O�#*� ��.~�Յ��O	@	 q!���c��
$9�B��j$;�!�y-2�6 �q�v��ue`�<�`��9���)��8x���^�}���=�^m�~�M�lp����}�`���b��yVe6ͅ��fN2��!�0v�TL�w�h�8mD���:D�]f2��!30f�D�>�:V�>��5#1Ewf��c:�b�ufY� ��]�3\,y�K%��R�A�	�_Y�U�Z�1�r]i�BJZ%j��*z�)U%�QKa�^��)
�p��"q����V�7�=
���zT�6�&�-j󟠎\�}�yOq;�	��^�Na+�RB��խx\ֆ�+( �9�ԌwZ�R4ob�_�*~k;�v�õ[І�}��K����Fh=�����#�_����=Վ#�d�V�>I�Hp������J "�?���MT=��_�� ���� �6SI�G���� �~����n�p�� ���! ]��wW���e#���>_�߈�� ��;�{�X+P��� ��w,F�D	8,A��R��(�eHtX�$�5H�_��r�8lB���:��2�(s?�
��8�Q��޷�C�=T���K�I�l�"�����C =C�-�~3afY�oZ��2��`��11l2�ք�v �mS�?j�E)b��h��I��1��0f�I D�lgL��D������&��d���6ٰ�,B~�	�P��K^�J�;\)�g��S �bZ� ��4/=V����)� �4H\�wIj(��b=��5���P��?!���>��rޡV@��f?CM�s�f=E]�k�����q��z��Q:C���V<Y	<]<YG	(o�;
@�fR��Nv vR
v3��0���"F�+��N��� |`�?;ڂ[����f>݊C'�p��O�C������G۰��{$���s���kH�/߁�O�s�F\r�j�7�N܉�֓� ���y��c@p�
1�rA�E����W=�6D�P�Ƣ��j_]�-�A��B!z���v�gìD�w�@"���|N�r^A�Q�x,�L7U
�a�vq݂��<���@z�||)�@!N�����@�	�Q��b�j�����eE�}��w-�~�l�Mb^�8X�X�:��"B�ȗI�����z��_�X9�?'�[Zl�w�� ̡�P��:ԅ��=���T��uTȻ��C���B�{�ɃV���eJ�2�;����ۨpW��&>Y��p��
qSq�(���N�9��>�F*N��G��)a��@N(	Sa�@5@��0�� �� ؗ Ύ`W��Ħm(6K��z)��#�j��W"�r=r�6"�v
�wb��!�w:�
���q'���\�C\�},��p��q?�M~ޓf�S@�P��z �S����V��������`H�Q5K��5Y��Ct1j$`�8����֘=�3��`�P����aF�0D�Oa1v�x��Zc��=&h`�V,��'b2`�y2&Yd@�2Vf�H=�MYu؞}�2��@�]̼���p4�!��=��'8�ǀTr��E�_�L�K|G����Ӝ��!�9~`����ߧ?��l�=�M�����p.��&_�O�u8�^�S�8�}?���ق;�P� W�Q*��n�s\[�7�������־�����O6�ǳMMxYт�[Z�f[��jŻݭx���m���bA+��`+�i����p��9ӆ�ߵ��w�8x����p
�s�I��ɩ�������������Ǔ��;#7��(ȅ��r\ـ���U	��@�6�a���f����6��Ip���dO0�U�ɐ/��|6�vl�?�sߢ�W�9��H"��D�+������p��l�"��6]�Ѕn����s ��������A���>D�
r�T�J���.�|�ߙ* ����{��"��P"�?V�.̚A�s��$L�|	�k�c͊��`�?��b�p�L �(z��6��g������؋�"���'�a�$j���F�����B. ����Q (����'�s�E�g���~�@�����Q����b�Y!���B,d�oQ�x�b,2+�H4[�d�2d��G��&X��R��Xiwk�N����z���m�}����p�+|�lE{C;ZZ��,�u��N����O���D����b� /�L�8���4C�j���h>���#�<��Ѱ��in3p&F�H�a�	04��4kL��qsb0N;a��b�4M��E���ǆ��j	�����n%,�W�ҡ֎�a���ka��N땔w��q=�É�8n`���~=��u�^w�2x��������0n�p�K��N
ܴ঵n���P⭓�@�4��gK���w]��+��)!�9���Kƪ�3X��#�g_Ħ�Jl-���K�`��G8��)�m��{��4C������{�Ȱ?w�	�N��܏�8�c�]lǑ���������l=-�hE��F$��*� ������zI��$�������� z���n��(�l��gDZ�w`��yJb��/��y��ȗ��O��`���c���"�M��3�?O�eb�sņ*�4��"�A�ݑ5z/䍮��'A����@\�&�"s���k�������RI(�<)��'uj�(#��1�>~�0��.ȟb�ԁ|}��ED��2����R�2��=��נS ��%@����'� ���ԅ�@. �KJw�O	����x�
u�/�\�E	W����,�<�|Ę�a�����N��#�8qF�)���H5Z�,�r�U��b+JmvbE`��lw����58p�(��(���CE�+}�@�t�q���:�~�?s��_� �� ��-�Ƶ��i7h�W�`T��ѕW����Y_����=�"S)
B &`��Q�2a:LMm��e��3�) �� �b��B�2M��4��@ڦ��u�w�����؆ ���މ �]�ٍ0߽��/A��� �� �H4��=�y���ُX�=���ܷ#Ƶ��MQ�o���Vc��*�r�R̷\��楴�R,�c�ՔB#P��7"+p3
�v�x�n,�ُ��G�.���~����ؒ}�sk���������!N�}��7��O���ܮw���6�¡F\9��G�Py��O7��x��R
�4����?܊�����f�U���~�a� x�K�/� _� �$�S���w�I��`��dץ(	؀e���#�lĲ@N7u�B6ߝ�A�;�u"A�#ۇ���
�ד#�+�Z�"��(�^�R���T,+��V��o-�|�e�� J���V�5���� ANy�$�� չ��Ť)n�$�Hq/V��ma'�J
��R�A�����=��/�]��Z҉|='��Mt+��~,�mS�-�w�� qxBEO�
@�Z=��@ݨA�m����u�G�B�~��0-�$@) ݑ)�u�6�EC�9�,Q�Y�6abDq7d�a�BD�R@bu�@��%H0X�d�H3*C��j�X�C�u����Z����#vy\������1·<AM�s<��-����[ژ�mh@���A1hP\O���Z�3_CH�؁�0z�$x����(�8�=��pz�u���5W1�����c��q1b4�5�ann]L��qa;g&��a�Q<&-�TؘbI��*}����\� �(V��c���]Ҭ�.�'��n܂��F�x܌�>�����
_�����^�&�d�$�Q��u�Oq-�1��I���Ñ�u�Oq��9n�yw���%��hi#�,���+��ru�u^oh��M��܎��v��Jq������(/�+ �� ����3 ڎ�c���M'�'��3�jŁu�w�;,N?w�B���%	� ��Խ����
	p����.�g�b���&K� !�t[����P�������4����?� �&�C=\ױ]�lQ�X/��2��X�	�b��L�O�>o/6El��۱=v�g�Ć�-X�K0O�+� ��Ԇ�@M@�R䍩x,��P��`GA�SڥHg@f2�_
�:�R���BR$��y9����>�T����}_��C�Y�}+��Z�TIV��� �$n�a �0�#}�@�`�L�M��=��S��!ݖ�uz��% �¥�pJ���j_E�CY���^ !�����r�$�緋 (�	D�[QH	�줋�@���B�y&"��kB��i��H���(=
�n�D�v6bur���x�B,6��"�x)��V ˲y��(�݆e�,ڜ�c��w��qǼnQ�⧰;��x�w�@�&��mG+s�������⊂=���	@?�% ,��K�0x*���X�]z	[3�b+�#˯�Ȓؑy��1�f`��Q7nM( �00��T����Q���Iq�fK�LlL����bqE�&\e�_]ªx��U�Z$����Fby��6T�jRK��M��e����p�t
a��5�|��T�EU�kT���_�:�9�s��Op���z�[����N�s�,x�E���wwY3�hã�v<]�X'� ���e���҆��m���-��aګ8@�j�C��a�r��&g��S�h��c�ѣ.�@Yx}�{��Ůo����3��*Џի/��l�TГ �PI��'������"��l����(┬����8��5��ۭچ���;����c���uX����θ}8��v/<�=�p<�4�$����XⳒF�M"�>C}�d�_u��u�/��cπ	4KB1U�%2ӭYnK�ҏ�t]҅�ubޥD-�0�r徕ȗw_���*2Ŷ��r?�Q�G�li���iE��2���� .�a�i� >�J��� �t��¿�G0�U��_@�^E�3߷Հ?��.�� ri�" ��_��@NX�Zd"�<!f�5IA�11LF�A2�������tDh�c�V�D�f�s���8�l,��A�Q>Q�� �l	�,�"�z5�l7��~'�8��j����vQ����ɀ��.��%���m�h��
�c�����]@�q���C��J�Oǈc1��n���Xx�/��~�q���S36�B0z�$�:
3gΆ��L��``ꄙ���~=+�5c1A/3� �}=~*d�]�z#�0\k��Q��U�5r��7��������|ݪf��Њ{[pwC3�����%��"NIח6r�7���z�k��Y��)z��yOq����������'�b�!��q��5��jĳ����^��ެmC}аxOh�n�fs+Z���}'�|?%���!>�.��d;����u����	N����'Ķ������}����"^\	�I1r[@�L $	� ��+�.���NH@W��$�Hv^�������:p�Ȫ�� �@l�6�����+!滭���>O-;�����ۯfЇ(XJ�y�S>g��5��:N�qk�۱�g=��+�c�N=����q"�;�8���;p$�*��b) �,>� ѝ�.�j����.�u�/!��h���UODu����v���cܖw�c���R�A��/E@K��J\
!|�,N;��EA&ɠ����6?G�؏ؿL �k����q����s�g��P��n�>��Pf5O��7��y�ۈA�
�˻
 �K\�H��$��@�\�@	U�
V�*�a���R(T�p�*>��-𻇾�,y����@>G=@�*��{��T`��4�� �d%!Ā�'"D7�:-¬	�C!��*9'�Z���I�|=ʀ~&��o����%H0-F�9�ز����(�چ%����q/�\����{l�����c|p������|��t=�eNЮ8$�*(����% �{a�W���6IƔA31t�pg ����c������}u0f�F��CFBW���Ѱ*�
]�Ph8a�TO����s�1Nw4���u.��.hD�T�7�B��S����+@�pmI'"�E��-{���ߣ��!�c�k�ۣ-�]�,�X�&C�Z��&ԟ���{���q~=j�Y�<���x���9�����z�Z
��=�q�+V��qc�}4�nAC��_��;ՈW[��\\X�#`-�v=?/��&��~n��C���Nd%�c�,�`g�I �����*�����m�+z��~��]��}�;��Ǣ�c�rf�������w�P\�_\�Ǔ���/�+�]�̅��#3'�,8�dv��4��,�� Q������ݬ���a
��,��
	�l�T�Q�-B_�"�%�s�؂P.���:�~Y�N�����@ʃvq_��ee���R�����*lV
1�~օlAyp���{��ǻ�¶`K�N�;�#���;�c�^K;�]���X! �f)�D��tU���K���sQ��`�L���#�-���^T�nː����}�GtT�ݑ`�V�K���涄!]�l�;ǉA-���
��Ϡ��k��CBJ;���*R!	�Rv�X q�t,�!WB]���� �{w� G��\���|��y�@�K'��ܿ�������L���{
|q�.����gVV�� ���-�^-�$Ԋ��(A�ʾ��W����<���.�~�	�~�T�`#
 ��`V�!zIf���P �$2�	ш�ㅔ��:I�ԥ�a�QbM�g���&و7��"�|$Z!٪��ːa��V�o�	�v۰�aV�F��l�}��q��6N���ŏ�r{=Z�mnlEK[=����BM��ٖ_�  ��k� L�ê~F�Q�p׍�/���4��iAfi6M���|�4
�����1�lcaSz:�!�6p��i���q�`�Nf�,@�{.t��.�J@]iW�<�������C�7�6�6��.n'���|��^݄Ƴ��l+jJX�7�.�����z�c4�lF%e@���f��<Ň��|.�~����x��5��?�!K�N�<-i��-x��/���z�����aS;Z�2�w2�E/����\t鷟��$��g:%����rqaq�b���qL\�p+vP �h@b�1���/tO���w����������";Yg��:�ӌ������Q��ak�$t-)�ҐuX�+B6H��ld�obHW��ἒἒ����\b�z�p�*��B����0"�\�k��������MX�K�)(�2|V	B9�����˶a9+���2�ElƆy;�+�0��Ey�v�݉|��6�c � ���
@�� š��oq|�!��Q�L�bdry �{��w��D�NP俔�� �v�$ę�V"�A�s�<?�?��*_\�K�s�S�;`Ы��� �"�JT"��/G�0+� �)���/����OB +� =~u���Z��������i<B�!�s�( ��s)	�z��T
@: ���d�Y���آ	��H�,A��R���@�E2-�!�j3E`;���F��!lp�[]/c�g�\ő�J����;ޢ�6E���,�Nףv�_� ��ྃ0��2
�����A�9��HvځT�]Hqޡ�����#ͱV%���0�`�HXTB�":�<��f`�F,�iGa�v,{n�� �iⱸ�Q���-��'�_�f��-�F �2�oץ���x�<<�������w��]�kٯ�����!Op�����y���Gx��^l
��\��8���n�<��째�����Y^3�4��������-�0nhGs�*(�!�쥠�$ �,��G)����D;~���~�ޣ��N�NHM:�@��'������8[+�*��Kt��ⶲVI0�� ���0L���XMr��t����B�4$p����r����X�$�%H`p$y,G��J��ˑ�
Y�e�	^���u(
[O�(ǲ���<r#�G��4|5r�J��CKw�C�u�����%b�i"�R��.3琎8�T�Z�Ko���v�X�@H�*Ef�*d�������8�{�6�p�	�>�2Jî�CX7w#2�ZQfI�6^�@6��0V�_�|_��ڐ�'�/������(Oٍm�����v���}X�
in9�d�%�+ $%�/PC�M�Z�����u��K	v�$DH��$:�#慄(�g�+QN-�큊@�*��#��r���
AGW�)�M�_�,$��X��DI���:���^V���9���Y����qьE�V,�u!\/s�e��h�4��k�7�@�4�=,r��"� �,�(B�E)�,�!�"�j��V�ȵ.G��F�X��J�cX��=����.�K8�p{=��ԂZ�e1�`�k|S��EOM0 ��������0h�Li,��Lwތ�=
�p>��l���/rL��7h2���`h���c =CL���|0n�<�Պ�t�N��o�����k�ˑ	�J�*ڥ[??�^�%��S�������7(u�-�]�
�ߵ�f�s���
/�1 op=�+��̾��[^���W�ʽ��{h8Ԅ[������������<��
��_���x����Ɲ��x���A	x��/�����Pކ��д���/�
(�C����CNs=E@�3��8�����~�0�wm����@#��!@�}^�/N����4�S���]�3�;Q �*�8�/�BVwn:!��Q��@�'��A�	��!�}�f�<� ����ִӨ��3Oac�I�O;�'�9�;����?�b�ylYy�W_ƞ�58��G*�����~�-�=|����m���$�,ކ�1��WcEp��Ē�2,�Z�i����ye��˱*e'���Ǟ�qzG�m�ā�8��
�e��wgq(�8����.co�	��8�d�DZ$�È��t,W}0��P�@���B$�|� (���
>G �E��b�~K�3�6g�E��uH��-ú�m؝+�E�g�tL�#���/E�H��$ Rȋ��ұyY��gv ��t��C�>$��a��A���A�9 �>���)X�v��� E�s��@#��4`��/FC<H{D�k����X,�͚ߙ��?#���V��q�]�p�xD&`.e"�bcƂ�b"a���|��و��E�e��+"��XhV�E�,\̗K=iˑi��[Ql�ˬa��1l�;�MN'����9��&�s��T�S�j]Я��^2�[�4��c�8oB��vJ�.�'���A(�V�c��� ����zI'�k�C{L����S=1vz�j�c��|$xm���W�̯G%�U�Z(5�]P��=��:n�dh^c�o@��6Ԯm�N�-i��r����,z���h`�_+y��̧�K����,����)#wps�#�y���ۨ˺��Y���yy�^�|�W������x��4X�f�3�-g+��jP���(�Y�o��(/,���8�v\�7�7����c��:F8���\.@�~�C��m�O~�݉�E&+|�<q��Y �YQ����?C�w�>�~��şb��i0�� ��nȉތ�'�6�V�DA�6��݂����l�A���/>K��K.`ӲK���ر���]���[8��.~:�U�_�Ǹp������l~�R�"� vdŦ�}ؑ��_���ؐ{[
�c����ݮk�t�.����g���'8���3��p8��<���GY�ö�#ؓwK�����(���e*�`�0T���V�:�������{	�����p�ǚE۰#���ȞH�(B�GR<�zQ��D���+ ��e��r�]����}(�z��������9�/m���"�e��D�k#�&��֙�Xe2�3:�g�v ��G0p��D\D����W�
V�I��~V�:���h.b���������O �3�@�)��� -
 �?T
���0X���	ҙ<b,O��<��<�o��..�B��b`|<���<q�2�|ĚbE δM
�ؤI�+�j�Y��3ۂ"�(�َR��Xjs�,N`��)l�:�����o���o ��y���������.
R8/��]v"ɵΆ�2h4F=�906u����5�U�8{���S"0fv(�̎A��I �潓$��T�W%����RO�8�_�j�a_'�"X�
oN7��z�s���g�}��9js�Mn^�y�G�^ �) /Q����7��0C|�s�����=AM�-�e���Gx�Ұ�ndݗ��.�6js� �õ쇸%$��RPڀ'�Z�b�fu�׷�Q�hG��@u= �P�RĠ�v?��S �g'[pj�s;ފ�\��%�P3vh�JA��1�{ ,8�}�W~!]�q�Z� ����!�����U|��k��� |=#������g���&��6 1x+�6��4l�R��Ev�,�l���a~	�
/c;�Y|{J��gy�����o���[�x�*ϐ��qf�=\[�C��*\�J~�Zq	�ˮ������8��NU\Ǚ�7q��m\9u���Õ3w�Ñ�8����cS�wؐq�Y��O9�u�Ǳ&q?V,؂�l��#i�o�x� a��-����T�������@���S}��-������r�G�s	_S,BN�2�*:���U�c�@��i%��%�9r��������*���*|-�;a��g���Te�'I��%v ƃ��J�D@�8����D���	����~V��Z�~V�R������33>3�ÏS���?@
��Y�P��7`�-�\�D��g��0���OG�u:汝�ϟ{��y�9�6���hC�l�MsmB��c������3��b��
$�F��:�mD��V��D��N�r��hǯk@��Я�@�7����7���\V(6��V��(�9��,K4fN6����0b�0
�.LM��SMO:b�X{⎑SC0vf f̌F��v\�}���b@�j ��|V���r��� �@�8<�Bh�zj��E�g�?݌';�a�����'�p���~� �-�,{%�俚WY�Wg�#wpg�S����4�Z�-\ϸ�[�wq3�6�����(� �$�)���&�N�3�ϡX��Ӣz����Z�oW@��f4mlA�V@�-P��CB�� .;֦�n�l��=/p��{�?ӊ=�[��p3v���s��$�/CB��E
�̓�M.|����?���{0���et�R������8Ӑ��%HcL������A�^�z�^}) }ѷW/�8��A�����|X�'�Q/	�q�6Z�H�4��.C��mX�IC���y籵�v�]E�(�/��:�YZ��+jp�����쾍�;n���k8�p?��r��J�2���6��Ɋ�8��6�������qh}-�n�ŉm��n���w'w���6J��8��&�#k�p��
���bo�e$9,E�nb,S�k�`�T�j�G!�K��Y���`= _�ߡBȥ'
���� ��J]��w_���� H��N�
�+�0�D������)~Y.K���,Ǝ��(�\�7�T"�_�2;���Г��'���B�
B)�*��.z"��#�Q�r��ub ����8�PU�wE�r����3P���D�/ă�5�{���TY�˃��"�_�	~R�,~f�Ŭ�U,�d��$+I�bd�ecV��	�g��1�u( ZD����+����d���pM��� PsE}>�tY���5�G��bD��4e�O)��Lf��'��i�e[4ߖ�$�6��LI�D[f!��i������0ɠPpjH8���Y����<�,�-�BݥX��I+)��c��f�.�;�?`��}�`D�	�k
F���ߎƸ�|�o,F��1��aT��6h���C��m Sc'hFl�,S_�:`�8+�턑�B0fZ �̌B��6���j�jr�q���������,�n�0�������w77���F<�S���?��'��L\A��mk���-��{���7���P:��+����b�\b�Wf<���{h8߄g�ޠ2�&����Z:+�ܻh8�����í��O�d�K<-�;ŏ(
wpK��<�ݼGxP�OJ_�ɲ<[EXی��h�܎�m@�.�y����		�D\�j�s���O�����c��{
@#�|���_#9�|
��/@  � ���'�n/��y:<���
W�B�w@[��2&�X`_G! _K�C���7}���0r�>�&���1J����H�݂�(	܀5�ؙpG
���*�C��*,�]��>eH�Y��J,�YͿ�:>^�$�'��!)��BW`q�
$��BJ�:$G���,Z����H\���՜r_��iR����GFD9��oD^�f&���Ȋ�@ւmș�Eq{p`�U\;�
5G�����R�m��n���+G6��B�/�� ��EHऎ�� d:3��^�ؓ{�a��-��ł��3��%ؑs �Q��f� �@��D^���W�.�U�@~�{�v݂_��5�|J zB�]�s�ʑ��~q/y�˻�UU��Y*|ԝ$×��1����C��X8|L"a�S)�ܖ����^{1����o6���\��g�/š���Т ��C�n,��Y���3Z�p�w.�W�y"�<����J?U"֖�σ�"VL)�X����m����7MG�I�b��P�T��]�-HC�V���D��Ü��,�B�,�[�$�U�.�߿�44p0��aG��d�~��,`gi��FcȀ�>h(�#Y����!C(á�e#g�ށ����6���qF=�#�S &a�p��T��§�ר�}��|R(z�s�@�K�>�jA�De!ÿ�M��[ێW��� ��C�x���3�k��+ ������f�W�
����\��E�q)�.g�CU�CTf>�s����!�(5iQ�q�9wqk�<��O����m��|�����K�6��Q$������{�]��K��ޒwx(�j��mx]���4
	���]"X\���w�f������y�vk����) �JxKx���C�f0�[��$ �i�&�p3N�����J�w �(�=@���`x�QНd��|��Ϳ��7�C�m��UC����5p��.~\z)1�a�/�=�ݙ�iǒ�p��]{<9�Ԟ7�h8�΅�~"	΃��`>��|�ypы��U?n\��unl܍!�eOK��y�L��p�k{��󋟅5�;pa�Uܻ|�.<���g�('r���}.��� ��E! y ���#���� 0��a�,�"I JB˔��� ���l�ڏҘ�� C^I�j��"�!��OS�:�m� �.�F��#?l ��m2���Y�
l��@>�b0�8��
}Q�'3��Ð������e�v`��AmV��1+xn�?�+v��( �_M�����P������Y��i0�����@�8�;j�0�E�0c�o��(+V�6��mř@~�t�9�����%��{���W�m:���HKq�a~f��(/<$%*�%P^�8�$��F"�5����p�t���D�����G�fɯI �a`�>��!��c��!4d ���F������=3�8��� !�1l�ph�1���#f�W@�$Z4N#GY`�� �S��U���0��}�_��~�ZJ@m�;�H���k��y$��!����&.�C1�^�7J��{���7�zA��C%�.���xA(��+SԤ�GM�]Ԓ����K{����C\K粌ۨɺ�jR���L�؀ڌ�����f�}�J�[q;��f?����xT�O��li^�l��5�m>�{���S)�{��ڰ����|����b��7�E��{�{D�����v�5�Hw �� �vy�ͅ/�o6X�� ��ØU���0�7#��;�ߝU�J��gWMw���{@_�6�l0m�5\�%�w��bo�����~��̫�YvV�FN�^X���jN�Ԡ��J�-�a�LO�\�x2�����p����(8�G�YH  g�(�W.w�$���b���΅��bL�0�
�a$Ł�kG�C+>�#��D�K�e��ʶ:�^yN9`!�pȯ.'���B]��*���}.!N�	v�/������� H��*ľ�c(Y�n�� ��
X2��^ԅ�_Bwp����"鎀�ъQ��j[̫��93DUt	}Y��<y�WCOg��� �� ��W���a�o���R�ޗu�w��}x1�Ux�Ç!��}��]y���B�=QH@'~|��E�5�>��<���6�^+>��3'>��5�~oV����g��a�k��_�A���q��.D8��������d�G3�c���������wx�S�H�S6�;
( $���h�b$�6��0�y!��3b�P\���u�&�C���Y�YfPbf,B��Ϡ̤��4�]0���ط/�|����>��?��ǠA������T��%#%5��^�1m:%`(�� M}
�54��B��zz�8J#��c�hoL���٨�bgz5�<��ܧ�������iO��q��k�W�SA)`���� )lG]ai$b=偕M�k����b�3���5"���:�a���Pr�i�q�����P�M� ���(\��F*%�� $�N �1��<���'x\�OK_���wx��/׶���6�onE��v�lkG�v��׎�+ocSy6o���]�}���������Ŏop���Q � ������e�
OC�~R'��n�妩�H"`H�-P+ }�ߎ��cLi	7���A8��:�^þ�?�t�E�N>������;H��K�(X��B?�1����)���$�,��K'
Δ G��p� p֋�2E�;����D@�;�eb>�����N.��0'�����ɾp��/60Z�����*�<ʈ�)+�d���R��`
֗	��w������)��@m�>! ҍ~�B �W �� ����Q,	���u�@Ⱥ�?�����g�2I>����B�K�* |}e��A~8��/��U��E7��	�������;r|�2|�L|�>- ��q{_�<C1��p{
���i�ʗ ޳9�`�ό���1��Ԗ���<��"�tB�Y�[R ,#�*�6 �Dۧ1�) �����ߙ����w���l�S��ʟa��0+V�,F���!�������ߋ6�/Ng)�'�3}f,��Y��.��[�3 ��^���_�W�=��������LHAfV*RR�����lm��p�0��#���##cL�����950p�1�a��#]1v��L�´I!��NC~�Q�;�Cٷp$��������8�w'��d�C�����%�<�w�O�}�3�@I��� �?���9��6��q���8�}��~ϰ�?�Ϊ/�ߥ��tJN�\%�p2�"a��Siq&�~H���R��l�U�O�$Wp>�
�	��q���S/����vWp��KU��Q���jT��@U�T�>@��'�Y�7ֽĝ��pg�k���'�����X��
�n�l��m۟`��ر�v�{CxMxIx*����D� x��I	��z���p���bt�I�w��ac����mQ��%� v����C�?�;��#5j,��zj�4X'����5�U���O�K>(>�1p�8�3���3�E�G�Q�r�I�$����:hE��p���q��Q$���a>����>��������do��
��Ɔo�#������l����ưg�q�࿇ 3�ա>��z �Y>�8PxEA+?:  ý[2�b����q����v�sW��h�.Ct�wň~E����{�$��X|�Y�3���/�������N�X�>V�*���I�!��c �}J�.絹L��Ԝ��1ެ��gE�oV�5��g�3��t�#Ȁ�g�>�f�1_(��53ǚ�o���OF�C�u	~V�.وs�A�K�BHOh*W0���m��N,<���c�|�Ϝ��N����(	�)|�S��L��Lc�1}ѯK ��A�Ɵ����/����[��ρ�g�	/?��fc��E��v���0l�H�0L�	��с��f{�H�S�����܆0�	c�8b`� ̜	]�5E�A7�`.\��Y��B-��I1<MJfK�k��fbV_���"�b	�ԜS�e0[�j���9�E� �K7����N���p�ŹN�O<�:S6S�H(\��p}ܧ��kz|�F�o2��Ӏi�p����!�LA��P�06J��"��y:�c�.���"{6Zn+�����Q���Y-�AI�q��|����j�U�o���-��m�S���;�S��փ�8U��c�t� V������c��c��@��" R��$��a�N	� 16@?�G����������P
�}8,�bK��L�����cw�!�9����;�0��;�(�RXi��~r �!��%]/�� ۣ�|�+���7]�ap$bjN)�`%
��|��{� .sЊ����^'����������4wXLr��T/��R���X�� �����\���w���1]m�:/�������^��+�Q��b���] �~w ��$! ��Y�+C]~72��n�J,����"�\.�\T�[��w2P$]�Q@A�
E� CYq J ��.	���� H��-�d����=!n���V � ?u�{���lܔg�% |^�X/GȄ�'�l)��ؾ��n�ň� �y�~� �t����� Y�������iϠg؉3w����G_H�@�3йL
u��8�P' �|��Q����u�m�K�?�m���K#
^�" �i��ա(����D���8�Y,D���[�c��b̵K@�=�����Őg��������w�%y\��yB H4�'����U@�R �D�6/=���|���=��`{4�L�W��mr4<�΃�T��4�L̒_� �~d�C����O|����޿W
��򃯷���?d� ���_q`&M�Scs�YCk����~��Q,t0x���è�.;����c�Ssf4̵�`���8��͸��2�������m��zw�xZ��O��R�Y,'�$|��Ǭ���ۨ�z�����]3nB f�3�c�45��?Γ�SBiw!4=��� �?r���Z��)�J�X�/�3��;#���i �!��P
@8������G�z��E�O��t�c!���BN�&�߉e	�P�zk��`C�ylYr;W�a��[ؿ�>V<����g�C�=@��X OG�?��ߎ��FƗ��E�ό�
�7���i�,�ǰ�O��\ ����, �@�?������XwGy�~TDņ��X������o�7c��}X0�V��"�!��G�CX��H��A�E�F����ݘ��a���R����ΐ"`�y�@XO�e5�Ϡ�+|;Q��w�� Bb�|
B4l4�a1�����#�'9�a�'<�B���a�4�ZA0e��)B�R�2�E�c�t�Uut� ~���b��T�a�o��)���\�8�#��χ��Q�T�Bo)2) ]�]F:?� �T<,C�a��移�qܟ�KĹ�"� �C �Aˑ&���n��>ó����^����  ��IDATp�b��)(�>{�����gO�<�A�B �٨�t ee�1�!xut	}5��m�>��#����my��ֲS����"���^Ɖ�f�{�g8+�}Y�K���P�y��Ǣ����ky��/�ߗU��+h�����MЊb�G�� �F�h� ���P�x�[-F�5�[V��I�b�G;� �)1Ι��������<�� (�v�F�C&"ĀQ�Y$J�2�1�w�Ip�f�0'
Nl[f��`����uRTBDO�$���������%����7��fa��q���G0��8! BCO� &���4N}��������@�o�0h�!���ȑv9�S&�Bo�\$zoƞ�Z���o�x�]�Ⱥ����q*�N�n�G���D���{�3y��C�s|���|�}�|�u�ut��9��p:�>N�����k8͊�TRN%_��2N&\ĩ��8�x�%]������㇤s��O||���%^�y"�縝�8�.$^����{9��V�J�E\I��+iWp)���jp%�:*o���.j�>@��g���5n�{�;pos=nkē]Mx��	O�7��Ar���c���ع��C y��_* čվ��T��.�L۱ި�>���G���Ɔ����{"�b{�n�\t�
`�	GV�VIX�Lp�E�G1�s���%N�q���#�A{.�L }<%�^��p����d/�O���`I l�O{M~A���̉&�8��0��;w�Ns��d'V��l�(n1�!N�����`�Ǹ.g�v?�8��,P|���P% �.��@��t���g����������Y���Q��?+�1�T@��K��"����^Q�
E����*X��zRV�^:m.WV�B |�>�X�Ϛ������Az14�� cV�b<�ق��]����d�
�?��ƪ>���ʟa떧��.�s�7�ZlfG* ��B�89�Y�(qaf	\��pa!�����e�$ _��`��_��l���q(��i(z�q���п� �4��g�P���M�7��^���m����3��&�ӡ(P�[`�8ghO
�҈C8�� ���Z�}����u�o%����1g4�&T�}@m�8���N\�G���dq*�|�ʴǸ���I��P���I�p�\N��+�*竒oszU)7�uTS�S�H�4_�|u\W�L�n��S���$��:.K�I�,�����7q��q�Bs+�d=���'����
_�q�[<]҈g˛�o�A�w@��v�.����7W�ێW{�c��j���	�{�㐋P6v}6B |) ��?' 	� >1��O��$	w�E=�7}) }���E���6�m|����
��X�+]Wc��Zl݆m��"�86�|a�0w2���K�;ެ�=u#��/�Fl��⸾4��_>=:��^_׏�>a=�f<`=3��O)Ф$���`7'vlL�Xa�͉��4?�M���4G�L���T'���d��1^�~�?�(���� 9e����_��aNy?K(�2�߅"�3�/�L}��J�T�W�T! "��!��8���4�=��E�[tL) b��� �ů��?�����a/-S�z�Y���R���Z �-_믇"�U���᯸n�j��j���	���1���4]�ʀ�z8�/ӗ�_}�t�`xzK����K[� o���q̟��=3
�W/V�>���tY��E#���2�啿�x�ڥ0�E�g0�31߅Ń��)�����P�E~V t�(���,B( ����81�N���<9B��_� |Æ�� ��_)�.z�t�?�G���`��I�2f��y�����_���S���?s�7s0�[md�a�L0n��Y8�qU�q-�)�g=Cm���w]��"�п�ߌq���zT����f.k�v�Q����G5�S������̧��\\�~����q>���~���R�=\J���IwY��ǥ���^��4�*S�L�A�M��i�J�mT���t��:����۸��nd��������7���v�sܧ�<�������,]:��
��64m� T m;�Ѽ�m{(��pe�m�_[�;�`q�N�:(�y�ρ?<?V~l�� ��d~R D����'���/�Y�S|�����_��|�3��ž��;v?6U`s�Vl������S��60k������N(�Ĉ��~����Y����͠���).�ȥkPZa����ɾ0�㉞��*PT�����n�\�Nᶓ�a>�V�~��9�����$���\�Oq��hG�@�(�6�cЧ1xـ+�I B�ս��f?�pq��źO��'B\�I ���n� �����z� ��3�Y�{p����`�z0X%� ݣi�b����3�-��9H��AfP!vEA�� ��}_��`s�N��_���K�B�Oq��b�x���:C��]�g7	�. �|-1@��6�G�M*%@uꝨ�Y����Y�B]E� ��������1]�	Ѝ��ST�
��BT�����c�
`��@� ���5����gx_�8	1�m(�u�[����Ǐ��K���!��^k>�4c�|xΉ�'��S�%����Hx������O;
�`�������b��"���D���?��I�R�g�����N�8� ��,$ L|^,�$�OJ�;�h80���v��!� �O�T��$�3��b�ׁ��/C�C _��|���(%��0��߇��E�?��7��^�����B ~;}�{
��q:����}( 1r�9Ə�A�U~J��ڴ��x���g��{���5+{����7ҩ}וu�[���oO��V\"X,+hD�tO����{��y��'x��N���;V�G����g��~���X�_`�)�..�����Gx���gVSj�ހZ��ӭ/���f�?�-?��������)*3�K B_��5�wm�MԐZq̀�;��u�2��F�C��z�;9Op7����z����V¢�~иh�4�jG��6\���WUa�֛ض�&m����8H. �C � ]V�:l8��co�$	�O
 S z�V� �� K�߅u�۰�oVy�a��z�؄��Ǳ=r��{�x�����l�#4�I ,4|`��K_X�`�S �f�S��B	p���\bN,'��b��Ƹ@g���< ֓���F��Ɠ�`9�6 ��v��J���/��a6���� �ժ��K��B^. ���t�������?�t� սi�K���Qk�"v=V.X���X��o��ĭ����%o�(Oڊ�)X���pX��"B�� �1� l�ݍ��ؠ�<��I���ś�f�&��߈U˱j�`=��[���1�����_$ ]���{	��Q�?u��^�"��@�e����:�/F����A �/�?��o����1b�2ȕx3���޺��u��CЎ����&�C��0�g�����`�{H��;�wN$������( ���3��0~�W���)�����F���8�z^����Ja	�K�nRW�'S�PȯT X��� �f��Ϳ���6��?��%c�5"��P�����������������Sơ��'R �R fa`/�g��C�0q�b-�����|/q5��P��ɐՕ�W�7�Q� QW��*^���6οG�@\@\���_�K�(|���>��v._r��n�z�m��ۀ�k_�bZ.�\å�븜̪������h9ۂ��W����\w#�6^Q
n��TrU%�x��1�O��v�]E�?%Bp�\Oa՟��ϸA�������nf��-q��q���������Q�<_�/V����v�[O���Ҏ�mx��;�^�ƍ��\Q�-[�!q�
 ;V�*�g��gA��� ~� �Fo
@���G��!�(��[��bG$�!h=6�n��y{q*�l�ۑV�b��0bI	p��OϦh��J�6��[
��V4��N�Q'&��'xC�+�;@{��F9Bo��V3��^#%�� �Q �&������KX����k�M���'ʆ3̧�B�{e�[;\) >�P6*����0�� ��B�{�`u����KXɗ 't%*�`O�1�(؏��۱9s;6��B9|}�v�e�M�,Q��k�*�&i3Ea#2���u�`���U~i�*>_�C�QTH��Ҷbc�vl����؅]��3� VGW ӝb�������t� ���@T�*z����v9��X b�a|�3��+���T1/	A� 0̥����^�4H�G[=�������[����"�=5b��wg�K��D�O���D�6� ��7��p�R�ϵI��*�?�����g��wL�t��J zv @%�/ QJ`�O� ������a����_� ��?��*~ ��wV��6�U�p���G��{#�'���?�'�@b�,z��8|��	��������������cHoM�V��`�0[,�.�9����G��~�����à�e�罕��@�UP��y���꾖��5����F���ʞ���%@�^:\P����������U�OP����z�s��ᐸ��\d�)�&�'բ��^z��;������V���ZԤ���=�pw�=\ɬAu��ʿ��>OP<�o�*E�*�:�S���ץ���"����۔�;����V���zD�N�3�/~�'��t�<]ׄ���в��?%��&l��	�~�QQq[6U"q�F�����<6����2��y�5�eØo�4�4@�^�� ]6
ċ�����a���Z���yp��~_�F�޽�uo!�( �����?��?��w,�Z�՞�9]�e>k�9����Ŀ&��a
+���Pk
�,��A��g��p��f�1�a=+V�����E+Y���톙�m0���Qv�3�ӇZb�q��J�~Nlf���#`��M��x��ua�[�r��-a3�ӽ(^0� �fH�)��a(�-(@&�p�D ����]��
�+b]�t�Q�����t� ���4�w�sd�bk�lJ݃�����^"�n&T�z�j��E�/.�+� G�����������*ŚX~v
�$�ɮ��Y
���OqhB~�~��; �_�����ß뭸�Zĺ���/A���߉bl��ז	�J,������E忀�q>��b��U�)��4�f�0� p*�3�ς��o�7d`�G(У`��Gw.�|La����K�顄{R��#Y�+�~�bП�L>��Q_n������E�a��c�����^",2�!R��'��s-��ǈ.�@?�]�=r;���2/ʀ�XO�G>��ID�� ���tȠ �P ��E ����0��z 4�lGl��æ�n�?ӏq����^�{���W�1����	C_%����s�z�5���P �1y�[�\&8��$ u� ��A X�w�� �6�E�O� q�_%���{���-�[�W��:������.�n���[^�R�5J@.�T�q��Zs5�u�?ҀʌjTR D����w+�S
jQ�t�p���SM�]�W� �+	R�
�� �d�3Sq(�v��+~��������x��oִ�qm�ljƹ��X�w��P 6\@��+ز�*�m�@j�( A� ($�C �2%���
@�^�H0�����2��P��Cv�"p#6GlE9���wcG�^d��ƴ�n�b؛�q���MeU��[{�f����	�<`<�&3�aL����QX��ܠ1Ė���-��f�3��)�c��{�0V�a0�
�i�Й��q�0�
kV�&�Ma<�����V( |�a&Ș_��.�.|t��P������� ,�Yà=���%ҽ���~R�;��:��)���-��B[�n�i�<(��,By�6lN߅46�b� _C��
�_. ��W� ?�y� 
�+u����K@Q����ɇ���m}u#�O0�F0�C ��k� q��c*ß ���U TSQ��W!�8/�N�J�) ��L ��S���9��>�a/�_�W�5�����o�+��t�z6�����AF�8�
	6%��_, ��B ����3�X�����P��5|N��V\,��ˬ��Ӟ�&�)*����W�ċ]�) ո�\�0�F����Y�si��n����g $_��m�pg�}-�sU�ץހ�{�^K�*���Г �%���q7��V�#�-z�GK��Ɋ<_ٌ�����PYvkRbU���>����ؼ�26o���1��Nec �<���� ��KȆ���b@���EЋЗ0�B8�_G`��s��T�e����q)����*��(s/�*�H�]	�h���	#�@���fz������pKh�v��x�Lt��4o����ޔ X��0�Ý�3��9C�0�hPfR4G9�|�/���Ĕ�73����8W�q��S��T�`1��#�`8�Z�,) �ȍ_�n��F�Q�p1��Y������uE�c�A>8QN�/����.�dO�)�b��� �����P��sH������,�3�$�3�?
� �~�S�[�"P�S]�G��߃ 0��*:{����H� _=!_& ����2�}^�)Z ���"��_\�/��/��Hk���bV�I���2���y��~U��n���/�������S >�~1�ۡ��ہ����W�%$@)�'�5�" ���o'���'c��a�W�1��F�7� Ѷ糺
@m�ˏ$@p+������������w-�.|�j�BM�;iZ����TjW=���H� ^M��Jr�!�p�S<����%�
��_�rJ5.�U���Gx��9.�U�*����x��1.S�=�$բ*�M�[p������R�E@! �̀��{����x��%/�+>��Z�|럣l�^,�ڃ���XUv
�ןÆ�a�E�G�S
�h�D�<&h��/�b ����	�T=	���# ����ߏ��P����l���X�["waux֒U~�"��~�1�4f1�gC�?��`��	��֘5�ڣ�;�zS��1�sf�BsZ Lg��a�Hl&�A�3(��^g�#&{�bF lg�qVl�=N5��b�8�p��h6�� 3��!�_o�t��Ӥd/(��~ "�蚎062�ueu���<�\�/t٩{=�z�����<3A蔁@G���C�[!R�B �Q��ś�>e�<� �� �tq/ uP3zB�|9����"�{��eؙ�  �ڨ9��o��>_�2�a���O��\:Ɵ������m]@��տ�S�+�-��a<<� /c����U!�7�?��G��(
�� Q���Q�Г x̙��W� �{iR 4) �?e� ��eտ�(V�Qv	�V
�|�L)�c���9X�] ��u���q�E�K6�3n���$����`?%��+ }�s8�|�a���oD�?F=�! �@��F����~�A����J�j�S���+����uo) ͨ)}�ʂ�*ӗ������Wҹ�W
��\�5\H��9Q�����M��[��IWq1��P[r��p�P��95�p��ҫq%�/���ݍ�q>�
.�^e�_�����zn_�ʴ븒,�p]� ���D@�t�dߥ <� <� <������mx�홧�W����(*݇��Naݺ�(/����	�j�P��Q0Ϣ d��Lq? ��� �� ���C����Q_�P��/��8m.�0a��'�L+6���3�0u�;���@w�7�Ca����5�Z�ȵF;B{�fs;�>�=����>�>�^Kπ5��Cn�?�zc�`���1�&��u�a15Ɣݙ����3�ͬ�b��)f6�� S�5�~�4��`K̡ H� ��F�����H"̥��^]�~O|�ݯ��� �u��(
��|�Z��ߏt_n��e���d1�O���V�u��B�|9�_C5���/[�[��"���?����\��S�,W����_�gP3 �H\�k�?T <( ☿�������? ���_t�w���E�/�1Y�ȏ\ ������%r��2Z:���׿��������������=��8#�Ѣ �c�@Ki��
@�}\�z���g_$ ��P N�qs��/pm��-e��X�˹��lK#������qy�5�c��x��W=�n�s!�����;� �����블X�R.���W�S����5<�x�ǻ��zy�?��/�p���u��J�j%�cġ�d*	��|J �~�S���̀OM,Gz�����v�O�a��5�@qް�`�((����vJ�_, ��o��A���`���b�W���xh�K�+�z�+L�{�`�'����cӉ�n�3�Lu��tO�k��#�0�!=�0��>g%`�7fi�`F0�f��cj(l�z�h�+̸ސտ����@?~9m�f��`D����t���1v�V:t���z�����	t(Z�,$H�Η� |� D��b	��~w�}O�} ;��U�~��߂�Rš>'å�|U8w����~�������W,
^E1�g=n=R�u�) �O Oq���
��
C�N8�� DI���� ��G�,F��D�8�|$ ���� ��w(z��������޿��o~7��|͠|Cz�FAJ@�ߌ��ǡ��&b��P fb��s0�[�dʰ� d������W�(\�}���N�fn���|1��$ ���ǋ�x���|@��&��o�u�������~��̻���^�G��F�`���\ǅ�+����P�k�7q��.%\A�JJ�U�_�r�}�=\���K�qX���y������*��"*+Q%Q���j�&נN��� R ��v�@2o�V�-ܣ�<.y�GB V��(+CF�*���Ef�V��姰f�O���(_{�����&����C�F!���_� �2�MT= l$� ���M����^Z�g��<��������7ߢ�7�,�o�������-�P��i4'�
�'�u��b]���XwN��pQ �'z�l��G;�|�7��2�GXB���g5>��㸯�^�qyh?X��oL
��h�r��$�s�tF�Ag�3���e����t"�cZ0�fE`�4?��vz��?����0k�4�B��)4�c� 3hQ ��p�"�j��: .i�\��% �(���N�����\%�gtG�veH�u$ļ4΀�c�"�9�y���" �
�ȩ~����y�{�aKE`�6,�ۈe��X6_���Kb֠$j�Dqd��9�X���2��d0�+.��}:*�p*A�s!r���d��]��*�|i�j,�^��1k�������2nV.؀Mi��'�*�� �K܇�?U�J |LK]��1~~T��u�ُ���8���mAϯ/�����@:�/�� -�7���t�t�_�y��@1P���hJ �ߘ!n4>�۞A.���N'^�,"��p����E�/*E�����G�d�
F�#��=�z�t�?�c���1U
q��X�v�{b=��ɐ��9U�w��	c�`@10���H�L�٥�3�� ����,�,̓�'�v�z�����$ }~?}�.	��~� �����&`��A����jcB?C$9��l��2���Ǭ�)�2��v��0�ň�|qn�;i*��6���U���Z�����C�r��Oq!�1.r?s��|�#�M��siwq.��&��YV�?2�?I���j��T�sIUJ*q�a.�/���,EAL�1�/rz!�Sk��X.�"�e���k�FW�o�*��JV�U��Q�u�r��v�#�*~�;+)=k��d�&,�[�����]�Ē��Xv%eg�r�9�Zw��_��y���������S!U��c&����|
�̢����
}� ��Z�U �B �)�ߒ޿������?�1�Rh�M��?�Ҡ]t��?��rq���F�fΛ%�]a�/��D7h����shr*�P"�0�簲כ�}N�� �r� 8Jw�3`�k����}q��D?XL��x@g�4�Ac"%b�Lf8�p��3����9�sX�k���`Si��L_�w�f�ʀ��A zFl/��;�I ��ʿW7�I((!Ι��/ q�=�S^�2�OځM{�1s6g�ǖ��ؖw;
���t{�s9/�|����|� ݡ �e�R
@����wag��X~�󕈁~[���"s6g��ƴ�(�4d{�~�� �������4�������U�n{�_$ �� I�� ��3��oJ�տ�1�H9�`.���J��}�)��%bP�;��A���xS��<P )A�B ��}�� �<�A�k�H) ���yV\귳�>���ݫ���* s) �� 
�?����3`�vKb��"��׿���>C ��d��4�jF����o�3#�.�b�-\͸��V�Q�����S\�yN^�W�5y��oq=���S8��*)�\_���A�B�b:e�bq��q6�.�.$�f�_�O��d��l�5��P��I�ązb��LL�����P���RR��c��e
�8-��8UP�Ք��L��*�ʇ�q#�ng��݂���n�=��cXCkM\���UXX�)K�!g�	�9�%/c))�xq�7��&6�d�w ���W� $���g�*I��a��}�� ���~������>�����!��٬�=��"�w�tq�`3q��8�
��h7L�g�!�0��!0ª}�Lǳ���(+r
��8G���#]�1ƅ����w�q��H�c�#�F�b�Hk��t��t�̹��X
�xohp~��O��bO�0L�Rc�`�� K�dJ	0��p�A�z �;+N�R����HD��ǈj_� �T ��L�����0u2�@g<�سi|\�)��i
�N��g�aw>�o	ßz� p�N|>ù"}/V��]�*ҹ�t7�q}qy�T6�i�<�\��;�]��b����S �	��,��3 �=4Xwqq%r]��b@B��� ����������S�(x�b�ӏ�/%�� ���S{n� x��tt����z���e��`��r�a&������=	�(����2��A zS �P�R �S �a*�P F���ؾz��%<��b]�aϬ�ɬZ�c�|1�.e�Ǖ��1����J!T�>c���}�Ky�g8���)�Y�S.P"Φ����������Y�g�~v��?.:��YJ�O��I�_t��� ^L���s8��Gi�"��c1U=� �<.	/ಊ��\!WIU�E�d^BM�eT.��CY��曃��<,LZ���r$��DΒ�(^�=J�^B��jR�5��^��d�`��_�tE@�N� �����8�S �ě�
����}�����߿����o&�^�!���9��P�/�b�����`g��d���5��`{���0o����hW)�g��a	���0�����`��?���K��.�֭�;��#����3��@k�3��zÌ��v��.�>�	�F�c�h�Mv��hM��4V�Sa�@3h�M0�B�9Д!]}Lq)�ti��8�Oݙ ?��S?�S"�_�8�_�|俜_" ☻+vq�;p-a�*��<׋���1xSI�h�"�+8&	@�c>�~�E@H@��.ؔ�+�#͉ۋ�D�V��)�/�#�=������Y ���Al7W=��@�"@~)����W�m���E�[w.���Q�V 4�J����l���D�A��\R��R �n�%����[
����
��~��� �z���q]������� � ��������C�<�{���~:�Jl�;Vs���7�x���ÚocqA�Z,�cB��f�a�kf����i��ڭ���2�Y��׼�o���W?~:��@.���8�Κ�Y1��(�f�w2CE���t�55X��L�/��q[��":И��Yᜒ�4`����P��� �)s�!(`1B������k���J!��;䔟��M�X��:�m��U�n"v�6x�1l���v�� � @j$�2h�0��^ #6F��6d�a�@Kx�|�������: ��m,4{��b���E�0x-�DlDA�z��.�뜹��I}�V����^0*�����\�!��%':�d��tq���mY��p�;�:#���30s�f���(��	%@{���Y��d��bl�X[�����Ɣ!f�2���b&�>�0�Z��8E"ܒ�6�"HCD��J^T��*�/!T�` 
�d�p�<��PJ�\�������z �u ���2���C {���$�,NI������J��}�W	��� ͑U<%@U<I�@mL݁���yq'�d:�~��?}9B �Ϙ�ߣ��߱���J& ��/zz/��Z�] T ��Lt��@�Jw��	P��m���x��W��,�����!/��(N�����/����u"(��'����������_<"�3�1�!�)����t��!/.�+���5���@\ �^\D-���i\�$ z�`?#X� ;J�ݔ ��/������~��~B :� ��,��$�=�O31��9�GcX�M`E7}�����l\0̧΃Ō��X���N��f5�ᨕ	G�,8�d�^7�ڙ��J���Xh��|�"�N�e�D��c����0��!^0��A��N��Ё����� ;����g���\fC���F�:1�؁�0�̇��b�+,�5��f���y�n�'�gxSP�(6�"�%"*8��x�z���@V�Q���%e����2�m��5�`�ֻ(�~��v�Ӟ�]6���2�ls�k�M!RT	��D��RLR�c�̪�E�K� ���6�� |K�!�>��{쳑�Pp�����}��ZC�ev��ſ�޺����l�!�!�0��� +
�4��a6~���+{����C[�g�=4�Xb�p3������4.�f��N�������6��ߒ`�iC�)��4�
����<��) S�sCL= |_�-�7����@�ti��/=�q��:ĵ䡯"�|� ���RHu/F
�4"����4���^�Lǥ��K��UJ8!	@�SR%	P�@ S�aY�j��8J��T|�Ń��] �( ��h�tJ O�h���*��?��ދ|��֩U��&@c �	�J� xP �] n�-n����
�F@2<���FD�]��O��6�_7
A� 
@��\�Ε��a������ �����Ϣ�U
 �[ ���^{]$@��$P��oHw��b ���fcL/-L�g���A��X���ğƾgq0�</���	�8�X��u8�|��o�T�-�L���iwpB�~�9=�|Ǹ�pb-�{�_��Ed�]pG���P��ƞ¡��qh�)������#��H�1�9.M��p~�q��cOp�$�)9>����x�I��=��qg$N,8��Opz'9j�)��?�3DL�[t?%�ƅ�p)�.\���*\ZyWW�C座���5�ߢv�;��~�����n�[�\{k�<@l�nx2 �� ��u� ���P�� ������AC�FC4�jx��c!���~� �� �� �F_ҟ0�?FB�k����;�!��6e.�G�B��qq�?G�J}����������l$��"�g�)`�V�D�A=��).�;������@�>��=X��}�B f��,��`V��i�0m�כc*`
�4�Bb2�3e�)�SɌA|�����s��(� ؑ�r48+x1�?�U��W�F<O\?@g@�[B�;�K@(�����=�<�E��U�c Ę i\��2`U�q?*2�0�K�� �� 	H�<mHކ��W!EZ�/!(	(��g8w���"�O��R f��g�G�e% ����6@�������"_��u���_�#��0�g��)�e��JSqj����-�B �d��|)�Ŕ��T�C_B��'����J�"@A����D���������8�O) �rg 8Ȣ ������u�N���)Y�S��(� P/ ��T
@���*���b��k��1��P���p�e�������1�E�k�+��[�����>D���oJ@��N`�O�@����@��}u1���U8�^�ү�l�-\̸�+�q5�tu�����}��\b�T�EUn=��p��s^�r�\�<���G8�}�����Z�s)�q!��/��s	|���
~\T�s�ɢ�8�p?P:~�0�[t	�(r��+��mĺ��(.����@����\H��%��j�5\���u��R�U\M�FerM�|O�i��˹���wq���-{��^���^߆����۝@�.�~��'�ڰvMVx���}�t�B(+� �|P:X�H�/�X9�W�0e��D:;@9��)Є���,�ρ��3���տ�n����3��[����0���;q��C\<T�L�28O��ɘ ���pghs��?�����F	������1����5��b:�A-*�Y�)�̤n����8�p��`�uV��}I�~2U<w�����ףxjP �Z!�UP��8���ǌ�;��;�3�"6s��S�ԅ��*��a���/�����%g��~yЊ�V!��SEh{a�q��2�s�/���:�6�is�N,�����@�����c����@܀H�0��!���I��.= ���J�E��z�y1 P���bx���g��U����" ��S����WT�#$@���;C\5����q���S�¥���(F���Q�B���� DZ�#�v��X�'��OA�K ��Mȥ ||�_E�w.�|(	��.tJ�j��1 ��KF�uE*���8
@\��9S`�g�|� ~]� ����8p��Z�Ӊš�s�!���~��}�z��<V�b��k\��ʢW����R�?G�>�(��;� ��^M	��O�	��b�~L��O�]���K8����A���P��X����!	g�����*�+N<��u)��S
�K��.|%�$V�2��Jb�zH�õ���UtwK���xT�O�6������a;�D	��ߎ�G�c[��l�#�<��Y��.F�۳�g���FVT�� ����@�
������,ަ��@�$ �: ��8c~3}��%sn_��Wo���Z$���mB8����h���c��`ro=L�/���b
�`J?V�|LT�Ҵ�qS�u OS2UZ�����2<�+���?>�y���>���8�f�-ff��V����3�f��b���c�gfֻ�]]RKn9���L�a]��������wߛx�I�xa�U�|M���[5���k8. 
k�H��-#D5 [� y3�f4�� �~ 4���K�obqѪa `�i����.� �t�W  ��u �1-��6�  D:��(��?������9����%�W���Ɍ2�O3~��E���G @�- �7�3 O�O�q��������{�?M�`� ������l�l�y��P�ƣh:�m2+� �����ϰk�e^�h���p�oq��oqt�5li=�~�C�	�É�Wp��8�*�a�1��U ����;�$v�;ƨ����)��Ǒ5�����_���J؎��m�m܉�Ρ��x�|��5|��5�}��/>��w���.jG�^l�߃{��� в;�肓8��N-�T��u_���	 � Wh�_���.�����־p+�r�>����O�
1��*+V+X���4X; J*]C�
 ���bt ��]�G���S�v_0^lGv�ƾ}�>w��މ���H~����P���3`��k����A3�d4�4�^9��X�.�"L��DS(��w��$j�=����Mb)���}������0=�V#3@ ���&@;���/ ��9�l����?F��?��m�J� ���ӏ8�n  2�O���g����L�R�[XT�r 4����h� ~�t�IS�} �Կn��-} J |�(Y�Ϟ�c)�֓i�I4�DF�b��4�xF�J4�x�􇑿��]�~��Oz��#ݧ@)ӯH��� �� �Hߪ?�&0��(�'����ѿ] ��t<��x�O����&F�[�dI^@�	���r�pF����"!�Slog�?�Sy�*���7�[s�i�{V\Įy����9����-μt�0�^w���5N��@3߉-��p|�YZq��	 ;�O����w.���c��g�G�?p����Bp؉.ihك���]�[q���8���2�(.?�/����^ ���k	����� �v5�S�;� �9�cN��8���B����k\|�*�٫����,��ѿ|�5�`�0��W���Qжq�ͬLM� �R� ]�$ sH�P��#Z�[� 4S�0����DYdb��1��o 2P ��;���P���.�n;���b8����~�Q�6)�O����K�����LI�?�4c��{PH�'�#<������mK�@��uD�ӭ���^�*&���דx����$nO���Vؘ9���F�_���~d� ��9�&B ʤq��k%M;Ff��z�`N�a�g�7ҍ  ���=��0 �a�jd�]:8�? �w���4o�}����ժL�)���s"X ^i~��x�ߥ�n����z@B8� ܄�����A���  ��
 ��%寉�?�om:�2}eſ�Qe�Y�и�i�I4r �� �d ��)N��J<�J ��|ߗF�H�u2x�,1�b�� ��Pۈ��f�+��,��W��6�o�� d��D�BĻ� �NJ�[M �M50z�� ����@�o6��  ����K { �s�l�s���[Xu��I����V�?K"�ø�.�/=��o<�޺��mډO_�������w�؊�8��$zh�[�	 ��U߇3�Ǿ������v�w����y�������i �	���@���Ö�}����8��aF?`�jе�a���Yqd.`�)�� �^� >��8��7xq�.,|��u�>��E~��Y#�� ��ed�jdE+M�R� �<4�2 Pk4"5��ը p�����}O�z"\����W��Ǳw���x�7�;��6�`�\ �q�	��4���Ǉ����7�3�� ��<hꄀ�Ӹ�и�Y���>����f<䇙���#�,�/���y����$�&�Z����y��}1�!�3�K�w|8������	|L �@�O	R#��NӒfi
�m�N�?�� э� F�a#h�CM �Z �&��g�C x����Yz ~fٶ�f ��~<Z�*����i�4	 ���[���{e���=�G�%��G4�=�b��	@���u�J�K������?k�� �;��	�
 ���������~���YGϬ @�%�}���N��)������>�΅W�����f��>���iޏκ����{�]��ŕ����n;��>�C�N1��N �E ؁��^�~���>���-�����;o+��{�_:�����H��~/οt��1�j�ߋ��ዿ~���j��6�? ��;��N��ҋ# ��
 $���G�g�h�����Ǽ��c��P��$�0���T �L�)b P�����h2
�`n�ɯ� �j ��ӟ0�c�Я���_;!��X��H�iF6���t_̾��|�<���߇q��q��IL�k#s�Iw���5�OR:1�w����1�ONx揎�������n�4���C��}T9��>�������i����,<5�~*��q������4���'��� l\+�
d�W!����F5�2�ߝ: d�t){&#��	 �6�����x��A h" 4G������w1;k�- �������������F�ޕ���J��R���Kw �	�2���d����)�������*�  @�gt� S���h�2	���a�OP�a#��� �n�h� ��Q�����!}�?��0 ��*��n�#5 �0�;��� ����h�{qAo�14c$����u�ilgd��濫����3\����;�������oq����j?��.����Z��]s[�a[�n��l! lŧ��{j���Z����;h����(�?���?pH�����+�4l�Ύ}���h�M8ك�?���/_��%Gy���VM�������O����]��@��݅m��=J;��c_`!`�i�Zq�V^5����/ ����ç�~��/]��E[ѲnZ�ۇ��b�ۧ���S(j|�1�0Ew��_?%�K@ �:4P�h�=0-�E�F	mBj��&& ЄX�d���1��]�@��?އ{~;�������|�o��ip��].p��.4h�1�~�DL���x�Wc1���w������xO��$��f<5�;��
�s�ԇh��`�#>ܦ�S��;<���*M}ԝr��ǽ0�� �x&�
�v(����=�Խnx�ng<A�x�z�����������֣|���xz�&>�ic��
���L% ���� ��K�rh>�� 7n�����ʞ��n�	phX�@@z<����5�4�a����i�?	 d( ��D���_JF�����P�ܡZ����ފ���h[���|McO���Z����Eh���s�u�� �^u���F��t h���ﾖ�}�C�/ �P@�`��o�m��N�����SA�/���YU�� H����2ُL�+��˂?f���?�ʵ*G��~��}��0� ��F�G��)�,���;w������4�\�K�Oez Ӌ ��ːD��� ��U(��!��p#J	 ���(K��ۘ�=�G����<��\B����Fab��Z���%3���OR�F����ǻ �)QC  ��M�7�U�$� �km��{o{ʪ!�=�� �  TX�����-���m `[�Y�%;�m��k�9�ZpG��^~�W]��ߡ��(v.:�˒h؍��}�ܧ��;�{�s�.\|�Z����S8��I�{���@��n܂O�r��@B ���_��n��>��(�>�)d?���st6���+�o����������M�Y4�Q�V��H�]��_:  N,% ��!��4 X�.���^�'_���ڄ�6�qu�VoG��}�����0
��D\L+R�	��tu�2Q����f	הFH��XYRi���&�i~�� qn��������?��]��{p���?����0�գx�������;�$�6��&��;�����=�۝�����1��1��0�Χ0���0�O�0u �0�aF�z`"�)�������{���S�ă3�4a`!`�0L$<�s�����G<x�3{��uƣ���G�����c�x� �����kN 4D:Z`�dW̊��
G�tG@����rbi�V��	h�g�� �A�� `dNÕ�uqX_���}u�����#硁Q}mTe����As
�E��O ��/ D ��o�m@�O�� P1 2ůY @�� � F����(��h��  �+O?! �-��#Mp�?Y���  # � B��:�,l �M1���o�� |��y� %{  �&;���4����O�A �u�Ylo��4��,����	;��c�``����k�E_�1��:�˯��4�.�ng�Nl��GW���ϰ��{e�����}��y+�k�Uӏ����rM�~z����D/�_�E��_�yF�W?���q���ػ�0:	=��'8\y�s^|
�U�����IV` �u���E'prٙa p� pm�78��x��ny���A�bV�K:1k�t��s_ڍ����h �&� ����u�"� m�6Xi��L�I3�l! 5�|��b��~����=������Sw܍���?���<�ݏ	��c����)����	��?����;���~����_c������C��]x���O��G1���4&�9	��0Si��$��+�S�Ƹ�r�����1�g�������
O�a��x�Q?<9����傇X>�k=<������z<�4ԏ��'�芰ifFD�@݋`	��%T�"���$ߓ�)p(0R2R@�dt�� (��(�Q @�ȶ���/����ES���nZL�� �Kע�ЁV��	혟��7���_D����A���&=�?��4P�H���#�_��2 ���ȏ�W�~=����ڹ�x����g�,@6�^��=)w��o ��,�+ m;��c��{��}�2�1�3���p�z���>]2�Ϟd8� ��6����wNŃ�s��| ��Ҭ1j?���#h:�--')��3��zA���K��?��w�%�]�r��{�\x�*z�ӈ�b��#��Ɨ8��"��;�}����?��u�Ը��ʝ�������b��C���8�� ��z		���=@��@���m؂��^��CgC?μt'�;������p��_����P������� �9� ���
 ά�l� \å��a`�>̩~�mϡn�Kh���g�,ڀ��}��� �*�#.����}�}E�d�aU�A �P� : � �a����F��qL¸��0�i�x����
����P0|���HHɶ?�h�~��"�A_>臠�� ?��G"�x4���A��1�|&��6>!�� ��h<�C�����@����;���c��z2����S�,���X�����}*��4!	�SL�C<Ʉ�	)�A�����s��A�+AFP	�Ū����,�! �}_24p4i  YMCMs�%Ѿ��@�d�_�k�Ef�5C�H �7C`Z��@����9�4 h�\���#ӁE�+�J�;x��]���:^�����kK^�{	"C�/�	  ��K&R�1}[� �r �W��ݶ@�w=�����0�'(yI۶�������G����_���@��/�zp�RZ�&�����}s�^� `�b�A�QV ���ŕ��gH�?��E��.D�_��e��E2P� �Y (MjW ��ۚ��(��� <���o �\
�3��5I�_< �d[�m�+��&a� <�{g��K@�߇� ��r�f���֋���o�}�k|��oq�/q��/���B_�	��W���6����p�+8��y�{]���*�GO�t :k{�{�>�y�,N�?��wasM7�+z�SهKN�R$  ��������U���=�s/^���/��Kg�g�!59P���L���h�CM :�u�����'�4��ګ8��*��=��k�R��-K�5hh|����m�,��6"�x%��xG0 ؓ��n��[b��V ��k[	H 5����禯��e����Z�9Y�1?{%f�ǒ��<�U��}�z�s_�^Ҕ�V�ՙVe���&�e��zkY�Q������&�y��]���&�Y�N_�Ui��XiY��5X����be�sX��iY�X���g���u��z	+�����ҟ�R���B�w>�=ۼ�*Ĺ�\s(�/k3�Ȧ ��f�#�);f�U|G×�GHV��!���& ]�:� @eM����P�/=��}4ƶ�1��ba�rF��ЖLc�l�q�{8?� �` �p ��- \��O H����K�?-���)m!��/����~#�q�/�~�<k�/Q���D�Y�;: d���,��,��Ѿe �g.L�7 z�_R���Y�  ��;P�Ъ  '�Q�Ll
�$ �;S � � 0����(�̯�i�7��- H`[�El�8�-mǱ������Y'�����Ϡ��4�u ]��u7T����m�܊�2Y�W �&_I���#�������f�_��TwY�*u��\���C_�.j7_�T�������;�����ܷ���.51�- lo؋��2�q�W���U�T����k?��zF���P[َ��٨�Z������x5/�~�[h^�>2r!.�ư:����h!�� ��6�#%���6L�O� �A F�2�a	�te��4c�u�+X�A���ͦ�g���,��~�z�}���+X��h�v:ϧ֤�^�^�ڴװ.��x-^m&����i�k2_�ߒ��2͞@���L�1˫Xcy��+��I>�J)�X�ԱW�z+�o��e,3����/`�I�
j��y,7R�#ͫ1����A 	��_�h=�Q�UYQ󬒑|_��� iq�;J|MЎ�� @��8 �T�:�[�����h��T��F ~�F���߳	�Z�/�'il[P �O��G#�C������~��5 �BZp,A<���%������ �"^+��Qnl3�#�VsPd! �1޽qη  c���}c~�8��+Yȇ&.R�|M�7@�h0p���3cn���MRK���4<�;'���jFٵ4����o��7���wR�ܧ���v���Nc�tl�6�`k#������S�9���C4�}���2�ߍ�Ru�v��lE_�t����i�%�/�~�},�J�dU>�-��+���y���<w��wa@M"�M%�_�S� Ɍ�*PKӯ�C��aW�l;�c����S8��"..��V^���yV
g�����PU֊�����[���e�(_��g���
23:\
SH� CX=��`" �"�G� ���Aj�8͔�d*3Z���&A�\���YX�H{���7��gͯ`=u]&�&/�:Q6�g��m1p�j5M{u��4h��-Zi��UbЃ�I�����<�g�`�#���i�b��V�ԗ�}����o9����\��:ϥ�xݥ��b������<V&?����,�<j�V���z�i$�~a�xC�����, �r��(s����F�ЕI�ʠYg��b�o�d2	��8�U��o+��e�O9�y�z����Vg]�מd�U�mF�����Z�'ffɌ}�Z�G���P��9�!0�s��k}=Ma4�PMa4�PM��N��9���.�C@�n!4�Dϣ��E+��&���tBԤ�/��a���X����> j� �?�ѿ��W��ki�5�����#ν�T��̣�` Y-�B3�1�Ҟ�*�q,"B ����L�@`:��� ���K ��D�wL��T�-&���US:� �C  � P`��"d���}K�r����4� B@H9����Zǌp�> b�2̯� `O#3 : d��M��V�X�<D��F�C�f�S,�R� �
��:�I��L �� � ��� �	J
 n� ���Mǃ�u��ߺ��T�WJ>�'-{�a�Atɢ@��b���#�o=�-�Ǳ���~#���2K �Ǜ����65�*���~6S�mo�ىM�[����F�����Z�����\5$Y�O׆������Wգ���oP��+�A�v�o��t�nGw�t7p�_7fmǮy��w��_}W����gq`�)t/ۂ99QQڀ��fT��������׌v��a�]��%��]�LS�&�\CH���0D��T�Yo`�/R&� �Q�U��-Ȉ⹌��B�(c=V��c��Y��2i�i"Fκ�3y��ږ�/�sWX(����*�V���s���g��9t-�g[n^g-E��9����V�
R	�����a�q�������"K��>� 1��H
�c�Ь�F�9D�L F�4,�=����l�peҸ2cx��D@%�Mzg�D�r�*�$���{i��+���,�$۔,�iⴕ��y�*~���'���?5R2�_���TT/%��~]h;�Xք��:�5T-�ky�6���}��D2|����І�vj6��
T#�@�@�����{�~) ��R_�WV�L򮡹Wk @ź�+ŹW��Zf@�d� ���7��X! W� �_�ѿ2�4���� xQ��GR])k� �V �  T��_  �  Re�! ���3��� C
�� t�'�����A���N���	����t�P ��7S��g���]��ޘ�L"y��Ւ.���E�򝍼��(^����(]�Ґ�(	^�R��� `>r�U������y6�f�C�+�b���#�9�e_g#C).���3���s4���"rҶ�$7��y�t�G�ȝ7�G!����,�x����e��*G&_g(�"ӻA%�I�BSF��栵d1��V`V�2�4����ō(/iAEq;�~1��[P�Ԉ��f�紡�x.��|�}yW �7r��lP5L!� �@*!��! -��� �ۆF���X�p?!�V���&��\��X��
��Wca��k�4m���eD�N���0��\���bi�m�d{��#��&������V�ϥd����',Nմȴ
M�_+1?�J^E���*�6����s��}�TS ����A��@ǰ!~��2X�Ybx �Q�L�N�Q'�E˛Qm����٨�5*�y�@Dռ?4�Q�~E3'T�E��l�kJJ�:b��[Pތ
�gyD�x��5�,������+��7h�U�'k�����-�,�u4�s�j�x]sQ;|o�/`"� :HF Σ��
�HS��|d8���g/ ��(ޗf�K��E�7�Zh�iT:^J&Oʃr'�/ z������W�9 d��X�� �S��&����yb <C�?��o7(�Q�F�6���t/�3�I���S�OSK���c�z㱇1�P�| SO�ԧM�>΂��-�1!3'f�iR&���������Ӟ2a�c)p| 3�D��0L�S������w�b��Θ|�5��A9`�Ӹߪۨ_M���4M�m��&�ھ}:�7��s��;�0��Θ�[W8��3~�w��<��/8��.��]�p���7�
���|&��I4��$���P�RK3�2g�"��b~3�:М5���`����G6�$��^5*Mu��be·�;��_9�I�����*a&�2�Ok�%�	i��ӣh*�� �"X�����䜍BO�k��p�H��{��(� f>ਫ਼,E^��R���at+��UD@���E0�ɶ�_��N��02�n+����ZD�2YJ��y����d[��&�尤x�D�<$�a��J��@�:d"fz&��QS��2jzbe�E�`��'� e�f��FV��Bi�a�n�	?+ �:6i�!�F���=��)=��� sd5��Y�� �r��o�,��Q,�/��΢X�CE�d �)��i��h�DQ�f~g���R��"f�	1S4E�(j�������p*tb2BdD���a�6���ӈ�i&*�����*v���2��]��~�h�J����/�s��gχѯ�? ��ժ�~ښ���_: J�_�V:Lq�Z[ ��|S�� �[ @̟�> |l )�� `t�� ��> ��)b`V�,��l�R���@��: dG� � �A�- �u�}K x�O�AF�7���@0F@�6F�6�ǚ���60��)x�wNx��x�n?�M�E��9Fu�`I�;X��>V�}�UbM�GXW�	֗|������W�!���
����c]�;X��&�e�>�myk�^��#�Jk-�c��봎�פ���l��"zk�^�J:���u�`}�kx6�u<��&�7Y����ų���ټ���/x��������-௭��ٝ�x^�҆���Lu��G��-�=��-��ԇ��=�P�	/�?���
��T�蟅>t��-s}��f.WS@Rͦ̡�]F�4�L�D6�>����H��HV2| ���&��M�Ք�G�!��� V,~�H
,AB@��sÈ"ƛ�wb��G{"�#Q��4�D�bE�3GФ�rH�'KBM�w½���2��,��H$�[�L�p�w&"�ȱH�l�yf!�=�n������|h,>i�&J��LOG�?F���5@��iP�5��$�F֊��j���dF*#��F��uI� %� ��f�F�OP�%�E��Ċ4� ��W��f����)ޗ��3\���b��GSQ��-�E�b�tf��D�u�M'�]FS1�i4nEO%(�R��lB��OH����?`A��rLG�s&�<[�\<a3�����#@�*m�}���H�.�9�N@�  �W��i%��B�� ���+h�e�e dF?�#X�ّ4��GL�j�>f�Sy��JS   �G:u���L>�2@�L�"d��l�H� l�.�=�C��_n�}��(1���e�� H �� FN>�
 b\
x�g}�z�f@:�� ��V��@���x�ȑZs�} x�7x�w��;o�����Z�_�~��r�G���v5�R�	�n>��M�45Ů�#�Y�e���ۋ�����V���Ʋl(�h���Xѣ����˻��m�u��9#������P�T�mwVmAW�L(�=�;�]-څ��=��I�B_��XЮ��o�[v'W�VK_{'�]Q� /����~���Uܷ�N-�������8��0B�QQ���ѯ{�u�Om�o�j�%�T�LH#d�7 ��Ռ�D��l�dRiH�4Y#�A5 �*KD2c�����2��M(1Ɍ��� S��V�OȉoS��D��*��R��LPѕ�c<79� ��!��I���Yх4B���!>�����H�,��@e�5��5ϡ	�2҈�/#�
�Ƈ<ĝr+A�k1ͭ1RI�r�^�|�ձR����P3�� ��ujn�7)5 e�ob�!�q���ʞ,��7�eI��H�{%��O2�d�C)~���
�r�jB�y��R=(�f�R��]�`p)D�3�{f.�g� nF6�l�9d#���$CCO�A%��Sx�yߚ�V"� fd%-31���3�(M�4�r����/���Iݛ��O�����*��&��2M�-b	Oq
�r	�+d6?Jf�3xfj��(��-�&��Sy���Pi!��0��s��M @&@oЛT3� H�����x�� �S���hg��- ��c ��H `I	 ��v:����,�S݃Κ��;�����k>���3h9��Y���*#NS���Mf	��Ⴒ�Paak�1�F�A�V�CoA�|;!`+E�&lV�-&ލ����ֆZ%ۢ�
hG���>�E�6� a�� �]�=�4���諡�S��{Ԅ@�ۨ��R���a_�!�wT<��N��'i���\���������_p��[�9�,�<g�y��}�6�­%A�~��e���V"�D\��R�V �a��K��ɇ ���ߢ�_7�AI_���X�e� _s_Vd3r#D-��1QI��.\���/�=%ZsW���;��h˓�!+��+^Cf�%~����u(��@AL;҃���pI�ע �Yq5��Z��UϢ:s>�
���2f�(���XYd��#/A�4j	�Ȍ�GC�*�C$�R�ȶq4�h�2D��#ʥ�-��m��e�J4�������4@?a �Ԧ3�? ңxm%��6�lM~����N�K�k���)v̲��֞����jp2����Z��5�� �5�l�ɷ�"�����d�,��<+�F��W�L�Iu��;�^�Y����w���%�%�hP�0�c�o�J 3��bf4o��>��P��+X�6���QF(�� ��h�������8~�"�����+rcY�n���rXGd����zdR���(�Q����S���҃ @�O��\y�+�%�& @f$| H�� �k�X Ȍ�; j�� Ĺj 03�� c0��{��=c1�wO &�;�`�2��hҠ�� ��0L�=��(x���e*`���t�j|\�}��1@#�ct�7��5�Ŏ��m?��k���Oq�ի8��E�Yx[ed ��J �;�v�:�>5��Nl�{ G֟����г'�Ҿ]���[w`���8�����G	;i��	[g�z [��&/F�*��^�h߃������M��ܡ�4������h�2Ж��޴�Vdy�փ��q��±%�qr�e�Yu�����~ͨ�[\X�έ�����˨%�h��p��v�ڊV����(!�'N�gD��x'�P��ʈ�7���xSKۖ�7�9��5i7-��UG�i�i6�0�0(��h�b�Yp�2iY��"[��}�M��ڜ�g���4�/���7Q�Ҍ%�/�>o�-�ºձ���h/]�
�yK�J,�}U��P�6�Q�3/-k���T�����V�
uyX�D���e+�T�Dm7�-FM�l�.EB+E�)���p=b��д�hPQ4��D�r�t�@��@ ��B��&{3"��k�w֤�G%#�U��`!��"f�"{�/�$��Θu��2��'��Z�䷷�\a�`" YR~UZFɛ��UfB�ų�^�H�,CKS�0���L�29�^�Y�D�����{��j�U����Ŀ������?���~#��`�*����I��o��+I[�{H�_�� ��v4��(7����]4��^�v�g��8�[.��sh���EeP�H& $���i�ɞ&��ҍѿ��j�T&�6LN���3��.YV����2��Oyi� ���]��"��#ϯD)�P� ��aU(��AqTJbP�t�� m����_�ҁҔ�(I���9(�' Hs�d9I@ d�� @�S�- � ����?�"˳�0: 9�|� fŧ~�����sWp����f��p�����#�������س���w�Ȫ3��/�w�Q��P�����zi�����`��}8��N=w_�-v��Q�3Ϟ#<� ${Pٍ�?��_<���~ =��	;pt�\|������a7����g�~�c�΢����:�=�`�-�` ί!��
V~�sK���Wpz�D�Ǳ4t>
y��M�G�S2��G!n�q3U9�"AҪVHt'��6���b-�ٟ�Zp����HB@)� �դ��uL�	�S���p� �3y��$P鄊��ȉ��ԡ�dM��k^D[�T3��-�e-��?G�_���<�V���"C;Z��bQ�(1�����Q�9���Q�!`5J�4�܅������"cR#���cݒw`��@����n�!3�1���}�Ө�hP���p�R`��Xa�dȔ,�"� F�z��72��w1 ��h���Ꮤ���`��@5@������ Ȅ+2�z��4V�& ������@ޣ����fB ?���0~]�, ��I'�I�^�dR�T=̔Q�;�f����]�3�0:~0 � [P �O,C~��(�Fqd�? 򤹓�dB�����"��^�t�E�- � L���l;��k����q��i�m2w� �a]� ���]��ӈ7�9�������	�`$�o�|��߰o�4���aϒ��a��_1:��[��%�/3�� N v,ه��.5���.�[xgןS��Ϟǎ��F�M�=�5g>������mܢ� d����-�߆S����˟��u;οy�PqI��@��j?��s��0?�� ��U� ���%�EWpl�)|��!�&d"B���ш2�S;���#K��. �_  �K )A�@ ��b���ZV�u�"��e�� S�Sz�@@3�J9����֧ C�O����7�^��dH�����`�1#�Tk?��F,m~��ܟ�H3�_ΩGJh9�UH�Q3��Ԩ�m��
$���x�VRR�c*Q[� I�%�(Aߛ�kH_��R@)����Z�� RiJ/jY4E�� ��}I������hn F��яz�{ `�I&����_�V�]� � 4��	 7F�.7  ' �,�@�d� �7xo��2Ĥ}ߞ~1 `�`�'!��o��u�{\�Z< $@�Nr�bݐA���-�L�wK���s�T*�\΄ 'B�!�'�m&@�� �<�@ �� �L ȍ�fL)V 0��a�( ��I��[ p�}w�C����e�_O�t�4lH�o��)��̠4���H�`2�9�n����}���~7���7G�15�ώ�s��rN��O�ƾ%�U g��6B��5p�mFی�Ͻp���1���/��=�٦ `���}e4��g�g�! �5=袁���[r��=�?O X@ �T� ����W.b��8���_z]U}����ݰ����6Ѽ߸��f�o���� �o�qY|'�]ĩ��W~���?'|E���W���oqz�U_�����Ρ��RP0.E�CQ0>	�#~��S�7-�,%��	Hvˇ����6!�����4���h ^�Rb�h�b���|HX�*���A��.yEI��Ǉ�6})�U����V4�Dc�*e��sQbX����*;�ׂ����&�e�B]�r�v/�JM�(ifV���N!�d���&4>�,V��*���U�/��_���y�Mn���5�)\���"�c��V�*s��R�7��Xٰ�iE��#�� DZ�lX@5�K;�t6`�!�ˡ��h�vd��G�h��I��HS�#�Ӥմ�v\�=�){����Bk��Q�q1�Sb ������ FGF�3h��� �����Vf]���G6f��4�� ޏ���~�a��  ����L��V�Vr���{W}\�JŨ?�Ez���]�(~��x�\��2 �x�4�L�����xg#�LHr"8	3ӆA� �@��k��I���S ]# ׯX�P `����Q���"��,�CA����t ���_��M!, P�С��: H�h-�_�$�b5JB���!��h�� � �ox���5�w�6O� LQ ���g��X�ga#�f `﬋��|Q��M�����f����`����j؁�k��˿|��޽�Ko]�1F�]��-�ř��<��U\��/?�_�T���& ���~�/װ��[����.��n =U[�W��5;�zv�݇�����9;���$ ���r3 pN `�W���pv�e]t�f��F�?>�τ��� QIc}�L�&g"nJ�f�q���Z @�]r5�,��7�����R,ma�| �B�)�du���ʖ��U2$.#����PfjEc�b�e,�WQjn����U��ha��<g�j�_���~�2����(7/ļj��6T�q��UF��j�궿���^b���<i����͟���^Af|-
��eh)]	Ch1���0�]@��	%�1��E4��DG��0FVaq�;��)� #3 )޵���� ����ЎA	 虁��� ����{[�K������u��	p 0Ҡu�2b7[ }0�/"`���B�Ou��� @��\�8h������!@��� �Մ�:B@!�i�oq�	�~@���wf�OE+�� �@ HtLE�LB�L�O [�f @�d����H��i@	��R@iB��� *� ��� �d,m@�I�QѼ#xOFȜ � �� ���Qe ���n ��w7\�@�q�^y
���9�Zw���b�������~;zZv��m�/܇K�~��<W:�~���;�Ζ>�6�@g����) 8��0�;�O�7aC�&\x�"���V��@�ջ�W��f�_�fmS@�W�K����8rS�K�p�U�Xz
�罅j�<OMD�3a4�`�=ዒ'|�|�'�L@��4���,��#vZ��,-03�$χ��@�G�$@�΁�&�,��DNІ^����$ �Ҁ�z��	K�^@N4��^�ݎE�bv�Z�h�/�P0�j=��6g!��We,@�y�˞# t(-�ƐJd��Ծ��Uk�E�/O��1M�1�a�
��B��B}�"tT��9�s�C|p!�C
��\����Bq�"w>Z��bY�ۼ�Z����
 2kZ"�L� ��5��@�p���m! ����j4m�0��A��*���,� J�tw�?M����ˑ�` ��r=]S!5���=���{ҷ���o��� 8R3	33�? d� D*�_�\�e
#kQ-5�$�%V�� Pº�(q�`�_��%�)#���I��QQ��yO����0��{	 a�T} h���@� ���Cme c�LM�ÿq�#t�c�@qp;6���@��Pw�	li>��Ͳ��)�ŕ��Ş姵� �N���>}�+^}}�� W�o�	��nt���ƪl���'U�س��J�o�ɟ^��~���⟨�� Pݍ3���b�'�\ՋM�"��k^z����� GV������]�=U���K h܅/>�}�;�z�wb���;��?�#K���r��8��2N���S�?Ǚ�4~��)8��@��g�P1>��"Q�T ʟ�B����XYOb*��dFo�޸���OH p�F��)޲<h	M���!�C��V����[��ժm��ۖ�Ƶ��8�k ��I�MlBS�rTe.@�e
��@�N���W!'���!#�	�y���g�Ն���(1,PS�𽖢u��_�<#M�Q@C�jd&4"�؊���Ȉo�!�
���y0EV#+�	�ja���*d�4* HOl$,4�$u�.�S�Hw�����Iɰ�X*��g! œF�]EH���s�[԰���.����H�
\'��¤9��x�0��U��2�����s���3z�u�0d�HshR��i6�Dfؓ�b�F�����a*e�����4�F�nHw% �|�N�����@̴lDN�B�t�l% ��G�>.�Ht�:�Y �O%R�,�r򞔎��MT��e������?I7�^I�%���]JT��#[g��K���.Ce�0��E3��/���D�d�$9K꟢�'M7!ف��`�o�F�O���+�]2 ���T��@A �@ �t�)�9@:����pa( �ƚhD	��҄Y(Kj
(g�2)5P@`���X	5l���FBv�m�D�,쩍 ��I ��E��T
����)4�t*!SS�Z 2k`�}aSҸ��� c� �Ʈ ��F `��E��4 (	jG#�-� �4��֦��FP���>��~�}��a��ؽ�4����7��@�at7 ���i�ݵ2�a�y/��v�܅O_����лpz�9�]x+�Yя^ ʻ��|�� �_~����_o�Vt�&*��k��c����fF_�v|�Ηj�aOϯf)�O �����ܭ�ن-� @P� �N��B `���s�Z�ή�W}�: ^q-a-���" $�j\*�
Cœ~���?��{��t4�'�#�hB��7d�T�2LpF��$	I��d�"V��n�h�:��U�	K�-�m�u����WGs��4����S�MH��T0`��qˌ�ΆUH	*��z$˃����%Sp-�XهT�Z�~RX9������%H���'%��>₊x#�P~�Z5�PZ<?CBR"*X��rF��4FD40	I� � `y Șt�k�Yڟ	 A�+f]z��H��i8�k1�K� Хe��0t]��_t�y av �j��m�fo�wd�we�wf��K��t)i��� ��: ��`�4��)P@C�oj�@������`���@ ��%J����'��  � # �@�ʪh��u�϶@&��{>��  I�2�]R(#����F�8�j�?C����.�1ph�`[f|���_�B>�jD ! ���`S�@@��Qn��2�� h���@�%k���N $��R���Q�xm� L������2x��Y2�
% �Q��u�p�� 1rM�� l��Ս ��?��4�� �� ��Fy��- p
[	 [ [�O��+�p���p��p���qt�4����4�8�HzW���!�������xx�q�uM���Ύ�4{F��jh� �+6��#��/q��+���U�W��:��{���̟����8Mp�1 ��w����詗����q���pb5��W4���Ҫ�q|�E<��
�B*P�mF����T3��~�5����QW$�ㄤ'�3��?ވh���*E�d� ����u$�Ko`�|V���gb��K���%ˊW��
��@�Y	Ӱ�BjU{Z:M�0�C��o-]���X��
*���h0��y,���6̩|�Y+���Tg�@�e1Z
�cv�<��PF �V,�xI�h�[�YU�h���[���|4W�T�B�on��jd&�bn㳨.��yM��T���P�@@9��h�ެ�%��o L>�*�, �@�	�qif�T�p���Gӿ4` >�k ��_�Z
�&�ߛ���I��Q�� @8@�C�H  Ne�C�~��QF� H���f5�OE���u 0 (�&�?@�� ,4��4@:�0
 ���Y�� ���P�g6�]ZM�EQT� �Ƿ�@��	�5d�� �����dP�뚂*Ժ)�v�ܵ��������Z���L�*Y=��Љ��cp��A����X��𩀇z��JL��P���d<���x���xJ  ��w`K��B�1�0�B�W3��B�qtW}���@��5S��������GO�n5og�6tU�d�L�K��T~E76��7Vta�����U֍�2m:��
���՛Us@wmKy�>p�uA^��`����z*�3�t�Ȕ��9ئ$ ��av�� �q`�	]vGW\ıU F�gV}���y��5W�Q�f4F��C��e3#P1! 5O���	O�?��G]`��ɏ� n��
���I��MNEo�Xްq��UF � +��8�B�vWjp!�M�x���Ŋ�[:~ie*���o����X+^V� ��W�� �j���E���%�Q�:�+ס�p�
W�1��5��d�2#;�+f��R�VcU��X��]��Hyh�\����X��<�	�k���Ud갨�%,i���F��
5EsPW"��k��ځXV&�  ���#�����HVf�vIڴ��d)+�R�
 �0��l�5 �٤2V���
z4���T�:�eP2����>��~�$�lz�	`5}]2��ڈԐFV�M�Eg�2 �31b�.?���f#���	 ���H�!��r���Wu�0�7��`�)P� i��%}T�S�/	 Z�� ����e ���[ס&�8�bB~�6��?�-Ok�'hs d�>O�nA���2�R�RI��d�8r��&�T�2�7:��77#Յ`�ٕ �,+�j �&}�7=5 �t����U&��4�"(�iFY�,B@+�٫fkg?���,@	�x���2��,YF^?яu�X7��6��o��Rk����!ǯY�����:>����W��-�$���_ ��m52�?$d���n3
�.(i�����Ӱ4���#����O`@2 ���V�h��?��)��y~�A������@W����E����3#}M4r��&�����|M�' l��J����q[@���)�wTS�U] M6  �j5��`[�n; p� p'W}���ӫ���u����[�2���y(�3��)
��Q3��O� �P��3w ��A�xeB% k� �A,�5v��7@A��IЉ�o�D�@��U�܊Yѳ�6_J�T�`�  �/�ieLm^b+Ծ���5h.Z��M��>w)�Rp߳�[�<�����7�C~�<M�͋T`Q�(6t +�A�ª�� ��H�_���%h(]�"���9(0K羅j����%X��2���RI�H# ԭFA$��6� �' � ��f @�� ��h�?; IO��Hi�i �F���O�� �D� )6 `���& Ց�� �j_�t�l@��\������M ����e ��: (���;�&?�m�L@�{�t5�_
��b���ob�/ ��D HR `t4X�|]��� @A����L����[XA�BaX�"�PL(�j@YL!� ��B�Z��. ���` $�o(C�o��W�� Ɏ٨�lD�6�u��`IU�5�2�	1�G%�4u �n� ��?9���8��|i�ݍ��[���{[񷜴�@)0P�� uG�W}�U��]�ܮ̿�|@��2F�4�Rn���K;��JK7Q�VmƦ2�Fj%ۄ��N=!�{����Y5���5��k�c{��i?�5�9[}	�V]���k�aߺ�XS��$޸R�D�"��*�XTOE�d4��$ wAʽ�Hz*��?Τ @e�5( P��l��? zZ:b2Û^�  T�3A��P-�k�(� �� Y��j��/�id�v�L)\G�Cnb3��Q>%�]h�Z��܀i���G�w5��Xȇ���ɨCH%���m8˨U&��s[=�C�<F-�Ê.�R-��Γł�h�BA��HД�W�8��� �4�#���6�ُf�O��6�� �ac��d ����t ��Ȩ֜g�I����H<�ߏM�@� â���n tI �![�
�,�- ҏ��� � ���� Q�g �w4�� ����P�<>����ôL@1�$���H �	4z[�W�؎�m�_}�i���
#��R�R����d $M ��3���&�	UP��kT��Qڌ���� �"&�� `,�^���5]o���> ��! x���x�.�/\�Ey�"���^�?�H�������5��5[�v+ަ��w���vU/ަA�M�~���N�Gx��x��/,���
����|o��7�ޢ�������7�Z�;x]�m���E������w�ߥ�Wz�z������7Kߣ�e	��~��������7���7���{�G�ᓖ����1��p+6/فO��Ħ�{��h�N�o~��ljo�"�F�2Ќj�x�8F��!Ӽ�0��O�"�~$?��	f z@ @�(� `��fB��t����	Hg���T6�s��JX��7� ���I�C��WK@%�j�@�x�"ly�2d�a�E:	�������J+ޫq����䶤1}e�Z	�A� ��D>�)|��նL�[A�gE�W�(y�/�Y��UQ�,CBlY$IV)ERp9U�DV$� @�  � T�� ���	Ʉ�,xC4X�f�4V�R�< �K�`+[�ڟn�?��/Ҷ	 ��*C�P�7 =rHi6J�:_��\�����{) �"\y �7+��`H�RWB ��4�,��TG�34~�C�  �h��B�Zz`G���Y�j&K�@�T�H І�j � J�O;���� � (� �M :�
 H��ρ �ir�4g��H�?�`o᳝��_�F��4{+ �d�( �D p�q'�G��@Ə >(}d���@��5�u}&���p�4�W jQ]�R5Q��(ІR� �������8F���^2�Fi��c=���I���% H�IF h P��:����<L�T�C�i��S�f��I�_ ��c���5��	���6��w���jh- �0��� ������������c���h"�2��48?��q𢼟��J�ד�x<f���Ip��#�<&N���1�w>p��3�p���.��+'8��)��Ĥ;0��i�����tL�m�Ur܉���y����q�f��yP��߰��~G�������������4w���no����c����$�Q�1���(HoGq�\��.@e�bT���9P�1ՆFT�U�:�5�Y��CZ73	N1Tj�S�ax�����h5~{�W#(�!��dMqSRϛ:a���ӐDH�C�̇#��G
�H�d�H��O��)I�Y[;;��D�"���?-��3�_��M��$�
 ��� �C$�*$�� �  ��&�R�����$^_`@  � % @3�6�8D<�$1�IA4~*%�FeU2ߛ�ϩ��~ 4����x7B#�D-�-�c����$���vX������$�����Yph�@&�a4�` ���Vx���|h����0����&�$+��N�'$���=���!Ϳ�~1�i<�4B�ٱ�3	�3�BH�I���8Y���#�0����J4mP!��&��$#��.���Z�³���ӷ\MI�-\�  =��0�3����W44�@� ����`.3Y��~�f ,�w'�)
T3�t�M�'�e��������z�#����h�V�Ɵ�l�I�U�&���j�j> 'M��� zԯds�����I��(@�@�o1
dt@@9��������ʔ�-j����6���:P���_�<�Gf�Lw^�T��
��?ѓ�DȌf='S����* # �Sxa� ��3t�&�(�- �c��QිpǓ4�q����i#*���!v��^@s�K���
��a��M�5��y�7X���5�3����/bN�s����Z̎[�ٱ+���̎\�������Y�E�Gk�\�F����j6�"��=rڣ(�|=���gN��:�y<��b`��B̍^�yы�0f�.ł��G�MX��)˱4u5��<�u�/๊��R��x�i�hٌ�gm�{m]�s[7>��<�����.�_���-y必�r^�^�sэh��jsF�X�`��E� .8$�;шX�в�@�6a�@@�8�B �ȇF�6��A2 ��hT5�
�EN865�0#f@j� @=��: �4�q��! H�K��F1|x�h�Q�4p>�1Ta ��')P3��`� �����{� 1�XV�q�4u%0�J��'y ##-� �YKE,�WQ� ���DҖ��I�߽_R|�4�Ot#X R�0�7:��)�@ a@�_dq*�! H� ~�~
 $��\5 02�W �N pO���Hã�[etN������G.! ����"B@1
	
��L����c� % 3���ڐۊ<��_�������2X{�˽%�X�u��[ `�Q��g���5�v�JLޞ��jh1  wjM �V� ����{"���kU��e76����Y��9�(�fCw�It��F�����m��l<�.Q�At������P�Wm����P�G�bCY�U=����m��e�	�q�|\>�O*t�sTtj��R�u}R�Y;�RFH? �`(�	�y�.nwV�H��ێΆm�ڸ������8��8�.=�c˯����j���ᬚ�*ά�tz�5�Zz��\���qv�	��sg����;1�n�oF�.H��@ϴk��a �T2 f\2bƧ � G ��hB�� +d��DVƶ� �R��
Xh�2�p:�:��-Y�̰zm���:��d�� @-I�y��W1��" T�
 ���*� =� �F~ ���%���'��H HG@��d��X�{�-��.�D��Ll ~F� տ��3e~ Ȱ��Yve;Z 3\�jR� v�!M6�t���o��%M6 �ެ,=4�Ot-&��Y��w,�� 0��u���W? ��j `r�i ,v �D H% X��2;�(�J_� �� ��Y��B@�g��Q�S�B�bh�	˚�p�2s`L#
c��f�E7#'�Y�2bI�+e�S>ϒ-�*�wS��[ `O�߇��>� 2� ��^[5�v� M�֯K�~]��OY!@:�:�� �������_���f����C�mІʜ 2p@fl=���c<~�Ǐ�O: �F_ϯ>�M�4ݪ4��XڇM%Z翍,7��c�z��m��u���Ҟ:�h�V�{l_w.4��Wz�S =��>�Vl�v��v���@�!l�{;��'q`�%^������~�����e:`�ŕ��²�pa�E��
���َ�85�8������Ѩp�A�N���ə4o3M<U3}�`U��
d�34�gh�O'!�d�s;~E(H $L& ��N�&��!0�21��I�*F�O��Hs@:! 3�FI�J�@sp-��d@��4 Т�5/�~4w�#`���!�	 q�@3��/% � ַT�zb eM��� C0!��C�?MLΗ�?%��'���$�^@:��.{��(-�])#t�u� ��� �"F��d;_�t�% u\V9�d�g�������T0d�H��'�,�@��T'B� �� yz>��J� 1�������~(ASW8�5��U9K%-sU��2Y�/ ��� ��w�@4�hWʹ�*�w'��e�/�?�޹�i�&�LM��BNE����9s������ ��'�����>�,@&r+��9���%�
��gm�B��PYM�p�:
��ـ�H�HV�+U��ĺ"�����  ���MK� J��M6���@��{������S��e�����-4�}4��4���o���'�����>�]�NbǢ���zׂ��m9��ƃ讧j��z߷��i�2V��G��Wc�k�Ii7�{���ߌ�2ܯ��>��>�D�2lp3#�^���ݥ[x�5�@Wc?foCw+�V�ey��m�"������ƽؿ�-?�㫏�ԺS8��y\z��0�?��k�~��y�[�]�ή!���V}��˯���
 ��9��s��@[����"P6�)��!a|4�'�G����:qO%#��$$�L�k)��G��	�-H�Ñ�E@ ��@�I5�	H�&2U���a���T��?�W:�U�����e~( H��ؠrD0��+A�1��@�}�ߚ��R�1����)�� #�d_�! �FoO�� `'��4"�o+۴��ȁ��u�J�K'��z~O�H�a��Y���'�#ѱ	3h*T���|B@>�CB �@���/28������
 �3/!�H�Mu�Q����j��"��H���t'�w$�LԿ 2�EH�v�@�G�<���C�E�w!�}�s�6aPaA@������
"j�Q�\�9�2ki��r��4��%�$�K%�$��n�� �V� �a�� r<k����2����c�a��C��gĿg�y|�����>����υw>���ǰ�q6�`75�Ew�~|��/�3k;6TӴ�����Ҷ�޽�O�����n��oĞ�{q|�Il*�~;��@�ƊM�TՉ]�����#���ʶ������8�+�����q�/�p�/_����n+�c+�\>��\��������-���-����y�sB�W8K8O8��kF�2' ���Ԋk8��2��;��sN�L��bZ���Q��Q�D �D��(��� ��c��<��� l�%�k��Z
,&S���&�_��PX9�>��̈́ �԰<d��@@%���_���f�b�2@�? H� 1ej��x�XA�[�_�wT� h"�AA %�&oO�4 P���� ����i ���?�]̟r)F��I�;0����� �DУ~�����o��{ ~�~. Hu��  M� �tM# �#�=� 09�y�%H��|�b�3(�_R��P��B@�V���*d0h���d����@7�[ `��	P3|I���  �p�mC���
���f'��cK�D��Y�f�y~����c`�q
��	�(��y��ً��;�k�1|��-<{��t��D���v|��N<{�U���o�؀�������W!�~��  ��u��؈Ko_��?�ߒ&�m�-ޅ�U[p����:o��=2Qm?N�p�Ǧ�-蟵{;�a�⃸�ug߸�����Z����pf��pn��qA���8��;F�_��B�򫸸��s81���(uJD�sJf����q��Ҭc+��	ѓh��	��ǧ z\2b'$���g�⟦�L@��J	�N|*q��	HoD�T$���S��iHbE��3�� ����0M>Bڲ̦f����-ٻ�^�j�,��3^���H/}��'��j�*��(�  �/J'H��B+\�ˈ_���r$P���&�p%Q����@�481N��|�4{%K��-�δ�d�@�>)���W�Kg��Њ� �3e��ĸl�����Q�$ؓ-�����d���Uf8�k��{l�%�� Z��4!����3��A�r�����܉ 0#� M�J���ɧZ�}��ʨ��!0� ΁�?=Q�29�F?U�?������F�3y��w�Sôx%�7��G�+��$�d	�+��}��N�����;�_)��_ �v �y �B@2й���b��Ժ
q�t�K ��Ĥӑ�lA���J��t2QM4�~��d�g��g�a�iT`&�	2+�48Yڰ@Y@����(p�,���`��������)�#T����2V���7E~($��>(�%�i�9A��f`�I�3 ��ޑLe�W��|�������f$�����/��ZX�U�7�&\���BMX+���gq3�f�b������`�(p ~ <�;�4aC�.��A �o<L�$ |��/>��C�n:���#������i�{�� p��ؾ�0.r��m g�<��]��=V ؈�k����Ǿ *�����z�u���Y����q��O10W`@�upSM�,9�3o]Ħ�-��r�Z�a��C���2ν�N������"H�?M�?����Z`�78��s�[��/�����oA3#�b�X;�h�7
�K �# �LNE�@��m@3�Q�i-� `!`�I�@�D>,26y��/�(�H��b�N�����)3U��u�K��YSq���` � �FI�^��)y� ��u� ��e� ]��B�`�`�y��Tt�B����@�� "��� �*�����m���V�S ��ê4~s�4hf"�O5ϼ�˕�3�%֑����s�$� 0;�S�e" x^�@��l�McdO ���� ��~> �o���!��-���ٞ�_�� N�Hr�C�sM:[E��u:M;c��J�L�#�2�Q  Ue(5'� ���X ��_iT �C��	���x��?��Wh��!��~v@�X_fJ�$A��g��U�O��VH�a�%  �? �QO�5�oG�R��!0i�L��L 0 \���e  u�N�Z�?1{����� �� S�z O��	E��4mYK h�͇�w�Y{��|�^����.b�dd����ك�����5l��B��������Ί> '_9��>\}��6n��j��}8��� @��R���9ASߋ�͝���5lj�%����.�}���9��Kb��C8��	\��Kl�s =�;������Yp7z= ���=K�L���pv�78��k�[�5�.�']����0���sG�k �gz!��я:��cEs�1 ��x<�H@ғ��d�� �;N2#��A0az�`�@���4V��Z�Ζ�.�R�/mɞ��o �j)��FR$�EЌd�?�%�%; �� C(=�FF�  M�����Y�R ȶQVM_#���6��m�1�O�4H��Ш&A��2ϼ;+�?%ff�/IS��R�m���r:!@�``H�<'�J��	S�;51��)� �,���oa������
 m! �hh" ��  �1�N�-���:�f�4�9Z�>#�2QF��4P�JJ��4#�@9F �u� �4�]��!�F������ō0b���.����Ń�4�*�CF�@�;�ߪ|�/ xI߀<����r�J��h?�J�)�ūfI�Q�$7Yr���?�!S�.�22�o}�,�&�BMR��?�%��H"@EL1��_�_ �? ��WT `���������K�	(H?��x��� ���b��}UU3@o�!4Co�AZw�~��r����_��m�'�Ww=5�Y�'^���+Nbc�Vl_��_:��Jm�w������`{�N��<6�n����?8h�R�J�@e'���}�M�]�X�	g�>���w�^N�~�N�|��οG_:��s��5 d���*p����3����[�� ���p~�78��*/;�?���n)����B��\G/d9x"j L��d@�D�Eb��@@�x�� �t H  $����J���JA2�:Z!@%`R}�'Yχ%�����^ҍ��d��ݝ��@ ��T! �C��V��x+� �	 � Q 1���<�
 R��3 b���� �hT{��g ��  ���[�H�T����@^ʬ�9��s�\��~�V
�vd;�#��eT�64PI^[����Y�Hz��@YiN J�#p��;��ym����13�U:?�Q}�B��,��	�J�K���$��� �?Z @� H ��u} �G @���oC���+-����Wi�o1�{���y?U?�������v!�D/m�8B�2 �v,D�c>b� y4��x&<�7 4{����_ ����h�R��(�5	�.dq���g�/ �N���U�/ƯIΕ2�Ɵ�I�3�
 ��K���	��|Mɶ쓾�^�dy!��G�WͿf�C&�G7�K.����c�2���^��o֘����m؊�����^|��ft�%X
)�������� �(M ڴ�C� Cҁ�
 ��v$ <�kG 6�:�V �;�����o9��?�v.?�M�{��i67�)�C?��ڋ�ƽ����dd�]�j���_�2���q���8��9F�]�=���8K�>�&M����@�f�fl��g^9��+6`c�F��v�&l��QۉS�C��8��8>��l���ke1��R��Z��@�1�[D �tg_�8�^k8��o��ά�g��|���>ņ�~�"�+�ޡ����P"�Ň�"sF�� ���� �H ��� 4�-$�3"A:ZG	��(>8�|��f�tc"A@_]PM��V�H����ߣ�{ >��4�ذj�J)��i��  t%�8� L"n벅�� �� ����2����"�!��s��N ɔU
�Y,��4�&�LX$�5��ۓL�k�A��D�b(�^i(���"]��,S�� \�$V�a�����'�"'�!zr:b��eT�+��tENbt��%tb*��(�`D �S?��'�5+SQ��T�X�D93b#�2z �g$�H���%���@C�E�nF���!`�w?�[�H��f?���G�~���M~M��$P��J�-��f5�� ���D08�ff��i�3�h�f� �D�O��D�I �9�N��V����v�I�"%F�"I�gR�4xi���� υ��,�Re#��@�{�d:a�|d��I�"����4SJ��$BP�#A��9��_�N����e�ֳ}[�ѳ��[�aG����5ĺ9�D 0[;�P�[ ���N ��Z��ކC�i>�/>�s�����k�0�f�^��zz�����S8�����]L ���?{D��/��) XN��w�t�=�8��	|���=7 t��j6Tn����݅���_щ��7���������0p������7˜]�⃯����� 0д�g�Ɓ >�! �Y�-N���	 ����N�6�����5�n�0����o>�^�� ��8��*��C" ؇ �u���8�P���O�R�$��Q����	q�E
�h�7 !��	���(Vpa#{��� =����4�
 ����C� ?�'���ܞn ��E9�������������R���y���<%A��8)�暩iR�i��4n�+���`�7��k����5�z:	^O%��*�'��(���W)aT���[�!�Ӽ���{՛���v[�����������T*e��M{�������.h(`k�#e���T��b�I?nk�F?�yFF  ��ǹW��Ժv@�63�3�2C  �
 ����-�4�������&�4k6@��e����3<s��"��� ���si�ل�G� �sY��]�d�<���-�F3M_��5R2|9���* �������rvw�Ŗ�m؆m}{��� ^\�
�]�T@�Da �?�, <Dc��Ix���,���&�AJ�?�_ `�{o# �a)������p��  ��m�  <��(�> 5��/+��@��k��7�}��Y����
:�����6�=g_���sҬ��U�Mu��k؂K�~��^lkہS�N㣲O�Ifo�ۈ������B��ݤJ]�zc�ft��������a�������=��K�aC]�����=���j���}/���%v�>�������7��,8�+|��^ŉU��5����/�@��~��������_���ϱ��X�Ҽs�KC�C��ʏ�Ҝ]��莐'�h�ш�l�����i�RN���K	 �b��g���J]:�I�����O&��T2RDO'#�FI��DV���H�iq| ��Y�
e"~F�Zf8Nt�K�u-d�R��b����h겈�8�\���ą !��!���@|�GC�xJF�����J�(sp_
��Rc0���h��͔��euC� ���@� ȴ�Hct��
:�� b�l+~��C�T���
���"i)%�/Q�|�.D~�b�.�z��h ����Pˈ����BF�y�D�����?!��G��51~�	�& ��1�*�<��A@�+�8|))}��|]�؊�G�e�o+�6����|-�|�x��⽥�AD���R�����^ @d�4�ۣH��'��e��p�s�fL4�o#ͿI� e�I�]2  ʅ @�r, ��3C �M��쐆4�T�Hh�)���h����J��� �7I�0����Fʄ䙄�  �  &Zǿ)��Cr�� @�O��"1���Aez�� y��<B@�h칄��~��l*��r��2]xOwͅE�=R&��yN�c&b��GM��O���|d=�p��TB�ʚ��ѵ��wcG�^���G��+�^A�s
�7��w%�n��p�#4�G	 ��� ��l@�? ���]��ß ��=6  S?���j�ƪ�<����4�=詗r?��$z�����}�e�^������Ϊ��Xև�2�����R�MM�S�����2I�� �;ͼ�q ����^��߭�K��T�5�zce�c����j��׼�e?/6Bd4@_�liڍ��]��~��ž�'qb�8��2N���S� ���i��g�7���;�]���8��
>�=���J$�Z�I�$���}`v���م�+��tdM1���L ��S�4�ɶH  � �H P�l ����O h�b�#�L HV `   � � �?��C�H#�Q�� (>��n�� H�&n Y�/�&D�'���ki�,C4 ���ą����=�*# ��� ������@�^-mL��%�e�� @P�! �����~���3�����	Y�h�B�0l
CV�0�������OP�I��}N+A��"VH�
B&e!����t�Ƨ�_ �+���5�^~��ȗ�	y?m���J4j{[d��I|�Mɏ��4��� ���.��EI�2@� j	 f�*>W�4�rD9�!�F 03� �i �0 ���%��d $�O��0�7:2�W �:��n X�f 4�)1�a �-柯$���@j� *׽ 9��i� 
l �ʠ�(�s6�?��1�I&1�d���h���h���DҎ:�8�:�#��Wa�����N���O�Ŏ�mxu�+��M
��u���M���� ��9E~�P�}�US�@��	pD��9�����=U��}��Msߥ&��)���5�N@gI�{�Y*S�v���:�Rf����>ݣH;G��Z6�,�΅��J��
� �N�23`g��V���܉~��Φ���~{;�����8��"N.��/��3+��������ܲ�pn��8��KZv	;��Di�F�ň������gz�f�@��<W� @$ J��
 :�P 0 왿�� �R �Y��,~^- Cn��6�o�G�D5��\c}��Os��d�BOtP"�GJ��-���˭��LH!�F|��a�HS��$P�� �,����˂ F?m�1}~, �S��ti:��h ���?t	��4rJ����K8��2Z/!�s������j1��	���� ���? �T�=�~����c���� {�/�|=��C%�o�i@
�1~Q���I��0��P�_��$��_ �3�-|/ ���6/��3��}��[�LM�ޔ,L�y�d]�à"ۚ�p�D��L�;f)�Qf���1�S?�L`&K��#��w�T���o�ć�? V6��ց]# `;^_��]�l�  H3�/ �����!�~���Q cX�Kÿ���q7u%�? &���jM�G ���������)m��5�+S�j���!TWͿz:+w�t�҄�js���b���d>F�e�xL��:� �B�������q9X��#������  �Vɂ@]���m����}��v�gžy�ph�9Y|ǖ^Ɖ�Wqr��,�d�5�.�{V����אA��Ch�	�^�u$y�"�ɗ�I�uA������Q�qS�%+P `5}[� �󟘾�왿(�M��?1������&+ ����X�d�f!�$�"=�	�� B�W�&�#�a�p�iȑ��$��i�4�@���� �$�T�{��k�d)�y]�-�J,���@
�� ��!�� ��h� �t ]4 �Q�P�<��\�?>���z'*C_�ɡ�1#�i���R��I6� �HS
oԏ �kGz����7���4�߷���%��|S�@s
��Y�k������_�� b������_  ©3	 3� @Fn���8 hJ���L� et���> )����F�(�+��M��	�2{�h���J�>� �\���� *[ ��!���a ���  ��ҭ ���B�RF")� ���C��� H�}[�	 ���b� xc��t ��� 5�0 s ��ccX�K������v]�9F ��Wy�d��$<��)x��7�1+�R��x�d�d������F�F�V�f�M�S��n�;%���v�_���z�z�z�wJ������w������Իe���}����6���N�x��/x����N��J�U~���n�Ǎ���҇M�[�ٱ]sv�o�,<�-����Q�,9��E�ѵ�>���*?��!:�����	 n�w	C�s )ߟ�7�	 1��{�	!�#65�7o2��d&&!��&�)�i e��/��������*���_��Q���q�G�O��'L���@�O$���0���HpL��g �%Ks�Ɋ*� �K �G4! �r�w	E��S~e�*��F `�F3�`4/ƮL��E���#i�Q�8!!�����\��d� �.8��5�i�)4=  `���� M�P�P��HE?d�f��'�s�h@�n�: d�t�  -P�� �ϡ�ٝ��Ǖ�_c��T,e���p:��)%
�& 'j�����ҏ� \/_��璂 ���3�d �����7>������e�ӟh���Ӎα5�������W�� z� T�O P��� Ȑ�i��4B�[�t����� ��h�"�L���f&0�gi b�b�I|�DF�#Y M2/�ə��B�W��)������4lO?����eğG�/@�_� d�!ۗ��S�\�b�xY��,B@&! �R�O�7S& F�� @��f���̈�F�� �m�{6V�������5���~�f���@K���w��/ ~X�� @ ��<�[L��7f��c��`"��&���d�<�o�������xx�����x��?�X��)%�{��u�?����� �����}�k,�ّσT|
��âM�����H�>���3ڎ���(��Y���A5(
kBid+*b:P�0�I�P;�sh -0ȼ����#�'�n�;�Fs�A�S("]B��hgOD�p��S: $#�  R @��	�!  ��0 �V2��ȿ�@�H�/ ��H�OtJC� h�qnY4Q�?Q��(~'Q^�T	�O6��p�R�YB�e�WJ`�f�He��"���R�	 a�e�9a<?\?F�R�\0 IV����b�:�R���$ ���f���x��>�������,5�@��A ya�P�T��+�^Dc�J�~����
�}�|�| �c_D�K3+�:$L+W!Y���V Ȥ�o�g$��`x�_��6ܔ��� �4w{�5|����#[C�!�#1�$O-�?2����� i �`���/�8
$ �1F�� `�����!�ΔM��p]��5��哏��ҩL��1���b��� Ǜ@� B������ѿ 4Ì4~>Y�D3�h������0��B&j�[ `�� �= �����A�
�����@0��d:�*����i��l��H�׈��`=r�@�xV#׳
�|_��
x��У�*E�1χ��(��/dY̛MSJx�i*F�	U:\4�QM�(���Dqp��+QR�j�V�8��1ͨKlG�qZ�і���Va^�:,�{�_���1��e�/xss^Qj�|mYϡ=k��W�ͼ���a^@u�u+!�Ѵ�����8!xJ$§�F���)i���&k���g�`�  �t�� 0>c��ѿabRx�'�o$Mc���dG3I�I��$>�	��H��'�a�#���a��  B �$/�͊�
��bU��� ��Q�_	��(�g�#�k�@��� ��IM>�fFɱB�Z5� � �}��H�+����un�: p�OM���u	�Q�
 ���ћ�Ϟl�I��A��L��e2T&@��/@~�b�/Ci�*TE����8���o����v�+���A�Xa���P����N&!��`t `o��F�@�������� ����'�o���� 5�*�V�G {F��f `4��M_����f��:Kk˷'�<%f�^��,���H�W�k��z��#R��	����@��(��L 0 ]t �(� �)��NIS ���f�� @�?��*A&��l�J��s��~Ȗ,�!�%Ou�Kw��� �J�72�O���4ݢ����L��~���� ��Zo ���I ��L x��e> 1��[ �G��W��>1�;�P��į��p"��z�����z��㿫v�Rg�nl���Y��k�bc� 6T�aCY/6�����.|\։O��,�Q��-����X��*6aSy�6ֿL�/C��K������/��������]���N�����TՃ5=�\Շ����m�@�Nlkك�m�y�b����3���;���O���380�ο��o��<��>�=g�g�q�w`��C�9�0vS{�sa���>F���i�&ǐl�J3#��r�XU*�7i�b� Jz�F��f�FJ�?�IMƧ�dzڈ�g���#LHA
�^;��a&I�)�Q:\h�|��p�{���X�L��A@�G�R�d�	T�p�~�M�
��E��P�@A \�V������HII�p����f�b�r;�А��?�&/J�����A�J�
�R�6��PuJF����� E��%���J�k�A�[ӻf_�G ��H� ���2�Q��Q+T�S�:\�}���K�>�v�w��"߳�[��!br��f 2� �P�PאI�	�7`1g����v�ѥ����{�^����ɾ��H��6�/�!��f�4n5�î����eۄc+�U�[�R�{J)���z$3pI"$���'�7�u��m�@��W=��:���,��V�H�
F�|K:���L>?J|�������gL� ��OsΣik `�1,Hu0P)T�d�=�ߙ�s,�qVɶ $����I� 2 ����T��U�d�a�3�I Ȣ�g+Y�1��U�o�t�#�g��%s����������3��Ip/B�+����;�z3y�2�1Se:������1�\���d�.���'�"l��	4~�dNQ*?ߺ�籥��Q o?�� �F�� ��6	�� ��x6�ml�q����@�̣�oP݄]]5��Y��*ex� 6�рK�����ۚ�K� �TL�[M�����/e�]b�4z]]�4y�6W �2@��e����=ս�죶������O-�M0�ݦ�nkً�� `w�a��{�������ph�E���9��;����٧�S��B��w�q�{4�( ��Ap���)��! ؃  T�5��@%S��4x�8�<��T����������T�5����S�P���B�ObğDzN��'z���A<略@ ��l �3�� Q�g¨P>�!��(�CM"�7��E0!��/��e�T3Cb�OPH`�D���"� =�}b��� � `b�n ������� "=�K0Hjؚ��4l��@C�hIy\�?>�8��_��v�x��c�Ǭc�NÙZ���2"�� ������p��_�Hb�����)�������_ ��{ �3���{&λ��K��i���=&������cܫ�Z����<$8�Ҩi�3�N��9�8#��o�e�A-��FS��p!�$"�%�*�N"$!��@2`(� Q.>��g�,�"d� �%�N��8f�43������FX'�NKE�4��ԅV��̟��� ҇� �G<����8�x�8�3�F��s�m�0��� �k>~��\��K#�F���[9�����f�:O����4}��L���{��Կ�hԝ������[ۏnF�h�ݵ�J�*	V�ɾ.YJ��k�C���u�����=�k�?���׬��s��������U;�s�a[+o��}Jj.��#4������9��s�`��s#���i�����j?C����Sj{o�Y���}�O`Ϝ��^�����L��O$���wZ<¦YL��B� �4DO1 ���4�*q�	ɓ�SF��ƉF�dO`���#Dhѿ��MC
#�d�2>�+IT�w.#�\Vh�
�/�3w �	 �"<
�:�T�V� �|�
	��D�aV�ق���������~J�A�I��,@ω�є�J$� �kY{>�KJM� �� `U�O�m�ن�H_��tI�/��O$�`Q�Jk  �#�����М�_�>��9.��� {?9���ב��iU����{�He �F�Қ �4�K�n߀E�,����ɖ�}҇`�m1��ɲ�??ǔt�:hJ���~��ʾ���g,�4���K ���5��j�E��c�h�C��"x�1M��VrN�G��� ��o
 f����'�4�4H�#�� �(�ޙ�)M�@��pMB�[",n���h��g�TB�� �+�&�I��������(�;P�>�W�� �- ��7��A&�@���看T+ H�/���S%�oҢ�Wᬻ�i�b���/n�t� @	 ���ŀ��t�� �n)�~[��������x��)x��v�ćU囹2�WC�lL�Fݵ�p�ū4��,`� �UmŅu�i����|N>w�����{Wߺ�k�_��%��R��V�ٗ�bs�D��j��;q��s�:kM�^���޿��>���v~��>�����,~�L�U��k���y���z
���@� ���ck�n|��W�ٱ�F~H���c�q�a�A�,��9��41��mb������ v����K��y�w��`v���b�`�W@"���wF2B��4]�� `�Q|c��@*%N�;E�a2�{>���ed�?(��y��F���`���	 ${�1��C���
^y� 㞋(�<DZA����ƨߕ �*��B� *}h��Q0@����H г q� ��~h��� ���� R��UE�K7}U��kR�e,���W �6`�k�ZX_f8'x.�B( (�\����ј��^�?�@���]�__���7�*��f� a2��e��M���0��毧���ݞ'�1+o*��+�Of�KAk�zD:��ZF�w |F�%�ʴa����N���Y7�A�e�;�߲����f4 ��7�g�HE��}巏���Kc���{�̽h愀�Q�A�(�j��ף�Q`F �  } � $��V�А�2>��B�71�7�@��2��wM@�;� ���;#�7���'�d�@ H �̪^�A�h������	b�z�.�-�J��W:��$�g2�,���/ �撧 @�:�az����g 4��!�@�J#Rݲ�l��a�����Ͽ���M1#bb
��  ��e6P� �i��M��{��	��m��j�;&c,!�	@�[>�܊n�����Ho  5�p���	ۇ5�Uoå�>U��;:v�«�]߫^˒�je'6Vmı�ᛏ�����y� Pӭt�K�9ga�}�1hd9��n��M��[�ȟQ����ˌ�-��l#!c���i��и}��c�m���k�3� ��.  p�Q���oo;C�8�m������0���wI_����Y�-:��;����4����-Ȅ�Q𙑂� >��`}(&�fB8� ����X�ǇT�@hH�C�L���
L��%+ f��D��e�B� $�7X	�����X�B�O�ɧ��3��4H�~�  �]	.��dᚇ0��s�Yq��`�CJ@&��� �+���*$"�*9G2���h��� �Yq�dA t�~ `��
�V��Bs �h ���C��� ��jk��� /�>y5.��� �w�ڹ/p��E�s�P�Y4'�C���M.g�Bp��u��������=�?�9o�& �2�ˑVO�Ʉ��d�J}U��P�4G��/����̂,ړ٤^ƷCV��F� T�?5�e����7#�#o�%�ٿ
 ���� b	 1�h@ JL�&)���  p$t; � � eƌ���Hs3Q��������5�� $�☄��C
e����zF T&@�6� ���`���� ��-C 5 �+K'�g�~J�EX7��sa���D�t�oD���b 9���d�2w���Էo�]�K ��S��ӑ�Y���w����_����( P�� z�w`s�d � �4�m������f3�.ُ���o���M�i����+6㓪8��!}�0>}�2v���b�/����5W:�zU��N�����M���ԥR�*���~[�k�>�x�N�s�WAW��t�$ |���bg�p �ݮevu��i���NcK�)l�d{�4�=�ݳOc��ز���x2c����#3���i3��3��� ��T�HE����
�"f���/��c-�,��iA"�d>(�����bdm��
]�|�u�(���t�s�.�;ɞ4o$��4�oM���H�D� 9����� �:�� *���� '�w&�(k� [R~�����!�]��Q�4�XV�m�b�,�O�� �Uz�/ P�m�4h@����H�|�`�fF�z@m�J\8z���?��oH 4��[.ዓ�����g��FQ�rDO�F��l�N��� ~� e����eh�\�V﫱,A�c��KԪ~�h�^�J�B��T��(X��},���m�`?��� �&#����������C�o-�xEz����oB4�p��{� 'B7�?�9�4��F��Hu��t	  �g2E��+���� R	 &7�?!���h��i���d*��o@�	l3*` 7�Ҽ
��S� ���X�w��V��R���^K�F�1���Կ����OQi��q)��b�� `Ti � �	e�����c��i<t�8���ѝ�p��De��	p� c����h�"�P�
x���̬W��U���V��w��ZSO���ډκm���kس� �-9�}����8��.���������;����#8���-9�}�]`�_Չc�����o��7�����6��;�s�F� �����UBI�kz�Y����O(���������6�'�!�I�繓<�E�e�23�433�,����V,�m��ĉٖ�Z��
-�13Ɖ�|�󪮞�ٞY�mY?|?�]M�Uu����|�3?�w=%������?�����{N�� �zتx x|�W�����׍��_r=���rv���̾�ߐ��S���y����۾/G����l����6I^b@�'$7�I�[d}i�T�t����^�'~(��0��?J!L�J��)df�C:c_3��
��6@@{w�6��-�-��` �h/ҡ>�N�A��^I���p�6b��	���gX�<���R�{� ��z��`��0�(�J��/�,�| �p�g�xU��+�"�2L���
�٦e� ���|-R>(��!IT�����D����G��`��i���i��t����i4�yo�����Ŧ_�Ri�c5�� �&�v�� ��8� ����)p��}2}����#;�����/���|q���K3�˿���l~D>4uXn����~I�ILW	t� �, `��:�g�e�^���:��v��#-Uc|o�&�ɮ����-��H���l�^�l���5��69���o��t*��/�� �2v�-���o�Ȩ��������ՆZyo ���vJ��#����w��$8�\����]��C����f�%\1)��	`x\B�c*� �,6
R���1��� 4b��@vki?���%����6��5_,���� h (�ed�j��-�\���HC~�4�" �o� ]FVS��@��>u�b�e�?�@O�_�YzIz�� |_͐����׎�q��=��\�Q>�*��!�c���_�1���J*���&��^O���\Ӻ��9:+� pf1 \��}��,Q��  �k ^U�_ \ �9 �� �2 +�����q%�o�� @� ��
d�k� t=��:����2�oK�_ud�y��~&Ͼ������!_��7����|�cߖ�|�grd�@���?��������
���mO[�����}�������1�g�ִ�kg������� �M��)9u��������� N �x����r
��郿 JΘ��L����=g1�����<v��� ��^��rz�r��g|CNݮ� �/�o���o�)NHN|P��m���C��~X
S����C�K��C���-��Ț�%X�AB(B!���K%y�J�Z�9�M-�)�֬Ym�C�>���
��������^:��/E:ͧN�YE��Q X 0U��E �  t��(�)�(�2�<��܍�ͷ�)�(n �xJ� ��+��+Th�bZq�  "UfA@=�C��j�HA�֥@5�ڊy�.��w�1|��[2  � l)4; �۽Sz1����e0  �, �H�_v%?(w$?*�%�]�5|J�J�l�Oٝ����?$�d��[	�#f6@�(�? <�vϴ��'����P^����=d�ѼfX�-���qN7��V�� 3�6����&�uM�K��S��� ���6v��/�� �1�¾F���� � �	 �  � s�1 �w( �  ���`ńm (�  � h Z�6H �Qa@Wu;jͪ�*��6��6�UZ  ��Z�>W�fԐ�nu.־EH��]4Mip���dC�z�= ��>��>꯲�ߘ?幛���l!�4 �$9�2������z�7� �G!{�B ����f	q?� FZ����#Z
 Ѝ�/� �#�R `����������O�\Ϟ�C3����	Dv>wF~���b�G��{�,_
�4}���?�+�M��3����|��_���}#?!�����o��>�#y О�������������O��Yp��x�>�my�}_$Θ��ϼ�+�} 8'g�=.���v\ �� ��|UN��� ��&gy���ߔG���|��g$��]��'eerD�5O��	Y�6�qBVWvI��C�T� ��`� b@"�JP�4�N�Լ���S u�&����OZ�K����w~R�v���^��ZࣝL���;j0�� m�7 0 a  ����o=&��0��`@jy�]��>�]�W����(F���d�CX � �����'� �  ���;Z?)_�{Z�|�Qy��g��g��/?�-�̾32�x7���3���5�U�� ���#�%/�iq3��غDn��w��7Za���-��I��f\���|V��� ���7���~ߩ��~	ٓ9���&f
g@����֫ )/� �|@�t֐�ִ]� � h Z��Qsi�4��7��k� � �Tn��r� dC�Κ �j'���m���l���A���~���V��a��s�@&�W�W�N󕘿�j ��E"k�$�Z'z���y����܂�[��o�{� \���Һ����f�N����h����~� o�� ��	��19:s!c����::�|��?������9<qZ���Ϟ���Ǐ��?{7Y���.o=&G&�k�
:��k����p��d����rb�)���~"�>�?��]O��9 N�=wۣ��/�P8c���9#' �;��/����} 8�>�Ⱦ���3{��{��_~���ާ1��3 ������=�o ���B������_��������ݲ>2-��dEӌ,o�*�[����9Y�2+�jz���,�,�O��X�/�� ��[�m�=�d�)ޣ��5��K#����J�k-Q�=��H{��p�β~�Ҷ�
��KƏڪP�F���
���kۿe�$��Ia����]�/��d�9d���>q��Km��B�+�`�t�T b)Q� PD97q4 Z �f� Z]��b4�����Z  �WH�h����� `7($\�@���3 [c�=������Y跿����7��������c����dg����_�<�_8�9
��^�:T.���9��1��^��h/�l)xط�3�b��즿������O�s;�փ9;��J���U��zv�u5 ��(����� `%J  �w]�K��h��V �
�U����9�^MƏ��Vb�d��e��D��X�*E�d�-�,Ɵ�"��5�h�z  � ��`�� ��KA�PiW  :+� ��r(���w���G�㢪S� D�`u�]= X} e��k ^� �V ��+ ��[��:��k_1 h-�B�[ߐk @�  � xtI 82��|�?�� �e��
���?#�����������>��ο�@���ߗ|�����<�W��Q��;�._�����)9������Q����+��=s�0��w
�� ?��8�����=''�O�΂���w���{���0���o?�g�A.�{Z~���&�'��wu p���<��>��������
 �ܴMnn�%7�:w��rS�a�d���a�C��7�����Jj��D��:^k Qj��-�CK) ����k�TJ:�7 �}%�j���M@�v� -�Q �.�� 0��� ��� ��7�]���  ^��B@�@������xhG�%d 瀀� ��Q!� g-��&��R�A  �v�� �5 ��� p� �w���.�u���_�N~�_����wr�S_��H_�niț�x.f������w6d:��IK�`~� ��)v�,}^n�y��;�����Q��i��/6�K)�񧵨�_��������/' ��>�m# �R	� � @[M'�0j��[�ۥ�
�'�o*��Q=�_WL����
y���i��[����+ g��l `DR��Y�:HV:�i��6��b�YݐXEbА6������^�� ��_
 �y�!���٬� ����96��O����2r���f�#�g�И5�ߑ��@�Q���r��''Oʩ]0����O�������<�W?\�l#���OϜ�3d�'gO�靧���˅����G���iSpB�Nk�@ �$��� '�t��)9����@ ��m(xϹ�O��]O�3w|U���<��9�`�<�
У{�f������w=/'w?/��P�讓��O˭��rklX�%��M���ֽ������rS�ny�{�b�.���|Xj� ��.0y�����%Z=$1���T�x���4��R����V��aCi�)�S �����Z ����R;������ �}0�PA��0)LޫƿCB��]�+.�� �Z^����73T�B�����%�t�Aŋ7�!� IP�A��F�@!@�5vm@s��4M����5c&wQ��ۦ������ �=�U��p�N�H�os�I0܉zܻ�ϻW6xo�;�e8x��G��ؽ������o��������o��W%w|Z�}�  �$HOI4gH� �u�W ^�c�9�Iz�ɫ׆���:M[��f�*���HW�����otq�y ����r�f��?U 0�� �*�(�=f\��}m����{�P�o���&_�"�B2}2��f�Yj� :�h�Ա�Z h�>G�D��V� � �� �j����K31��a�j���1���J @`u�k � \�z�N����xlM�#����L���#d���Q��2�G�::�㴎 ��ȶ'N�����5���GF��Qt�Ǻ.�>?l�	�މ|�I91�q��|1q �d�
:k�� �<�N���S��I�?w�43�zN��H  ���٣[��љ�� p�Ϝ��(Y�Sr~��ra�s��s�sr�?���#�?���_�_��rj;����=H��L�e���A�1>&7�����;��}����������F���cRU�UŨQuň�*G���ՃU
L+���cG	���t<���n�!q As�4�d��fh��, ����*�IT&�G 6�ג�c������� ;����`m������`�!N�ʻ� mWM�ڵi�~�,�A�|̭`@�(P�	�G��6�E��F�b�#�J" �JQ�:T��a�Hk �` �@S ��=��YK������U6 $ܳfLx�ߐ ]��V�r�h�����'��d0x��F���}�5�vy���E~�{��/~+�?�lK}P���`�$�~�10�vI �9�^�p�-�:8M_g����~�jۨ5�Wa��}6e5�K�O t������  �_�� @\�� �� �� �@;[j����|�t��s% ��+��vi,k�TWBf_܎���v3�X"�M��|
%M��UuJ� �s. ��& ��X�--�ԧ��*�6S�d1���^�� �;2�?��9�~1 ���T����4 |���	T( ��~ ���|_۫ ���Zy� ����f�3 ����-oXatϯ���i-0}������F��k^�R��;���k�MoX/�[��[>+��\����rb⬜����:�~�	�[����O�����ʉ��������:5|\N���3�'�Ύ������i���|�����,!2�ӋtJa��:>�� g��;��w?.O�}R���eyrϳ�z|���8�z�Ǐ�~V.�=/�>l<+��?/��>.+Jzey�F��3(7�'��Ĭ��~�\߲O��C��u7 p���=)�|EŘTVN�5.UU�R��0-�j �
���k&	4wMH�m�V��5 �դ0�c�+65Ul2s������������i�� ���C�aiC���3,�^���
 j��@F�\��1c
�N)k�?F�V�g�U�������}����u��D:�V�p�	�NE
��m)���N�R�Fίf�͜��*̿j�R5� ��k��������>KvM��^K`�qޯ�蔰�&L@@W�k��U�� �9x��D�;e,v@��I @�_���������%��~X��8k7�,�  �*��K�}6���ke�l6C^ ��k�[���2�]ۡk8���N�Ku��&��;��� �����=R�R@@H( �8S @Q�w��R�_�+�@�0��-�QZӵI�J���/ ���lwR���;�ɘ�4��a��~q�$
;1�K�K�d֪�D�u���s�a��dč���4�f���$cf��|L� �w���?�0�v�>���1�G�s��1�0~���2~[�9 �l��|�ġ��2tVA>\���� : x��V�5�瀀뀀�_�Vn���%.���_>3�|f��|i��<<��<�@M�'�����"�G���#��dtpT�[���<2�E94�%yd����ė����E��/��?htt�Crl�a9����9K��㳏ȉ�iͰo��N=$�'����!9��9��}TN�=.g�����@��srb�y9����{N�=+��<+Ν���:#wo���h����-��r�{������g���v�A��N����{�  ����x^�aUa�ծq�`�~   �x��b�� R<NՌaΣHg�ðQc� &7H����Dƿ�d��� -:���� 8h �����Ƀ2��4��t ��C�t~x�X�ۙ1
�S6 �MM@�xs� ��. ^�%@��	@ 	�J�� �RW1*� P�X5A�4�cK���:Ω*hu�N�b&{���^Kj��l��~�.D����Z m
���@@��3�P�n���KFCwȹO=%����C�:+ӱwP�Ic��1��d�&���7���m�
dK�	�WS����e �R��r ��X �!@`1� �@�&I��!`ЗV/�~'�0�/%�G��'���Cc:�h^�$�R��?�� �6L��� ���o���n����&+ש~5�_��m�x �������MW Ξ�N���-�n����ɛе�[.o~�J��o����u�_++��Tʯ������nL��z���Aܷ6�ǨY<�ئ彵Q|�ۛ��{m�t��[��_�� 
�HIhe��W�s��	�udKu�z��4H"�QyMPo�C�鰗d����n�&�ȚF	���h���1)`�x{̀t�!wTo��i%n�1֔v�+%H��I%��³|MJnΫ�*��>�����%:%o����4햛�ȍd�o�W��O���H�TS6�  * �J �
 �uM��]S`��#�yH�ƀ�QD��¬]Ze?j���f̻��WhFM�~[-����洚j��n�Jw�������Z���2 `g��5��V/���y�'�kS@n? ��o�(P@�[�	�߼@��-�k # $R�#6$VA&�J  ��Q`�R�b������8ǩj�Ⱥ9�:ǻ�򦊩<�Fj��l�Wū�%Y5�w��j+�qVZ��v׬tb:)P�g��%p���.��;����=�m���n�/�CVL�p7�(]��[������Z8
�b P���-)'�5�k�B��[2C��r�_��}��Zh��e���G �Q �X�ךz9����S/ .U��V��@��l"���������a�(Y�ѣ�#~E�0�\]L�C�l���Z; E��{9 �_;���T����3����	5p�_�<��������S/ �j ����p�?�M�Jf��W�U�^&o~=据�`��  ��IDAT���<�&�7�����F a�x��b�o�;@]��Co6�:�`����$tK����"�˻�a%�GӼ������ֲ~�����!��x�]���FE��2�2�n�NW7M77Q$ك���J_a���Ɇ�~(� )(d��6:�W��,<����(X*]������Ǜ�r�1�1ϤL��e�7�vF��[e<�m����M�9�����0�� �`d��b�I}�����Ni�x��w}H��>*ɾ�Ie��喾wɛ7�C����U�R]6!el-��1)'���8\�>�?�<��ô0�Z�^���{0��tn�5��	o������) ��� �5 `�1;�����Um-  �k��W Ц 5��� �^_�Hk�����
�BZ �����С���!���-P�b\���=� ��R5d�(�yM  �����EUn��m��o� X �"�ס���j�< �Z � hg�M��e��l��/�sN޹�?d��4�NJCޤ�s���)�u�WӦ�f��� ��� T�j��]Z�oIg���ܿP�Z��YZ�f�M:r��U��ʵ�Š����t% `�h
�F� �['� `C���� �sd `�" �rǸ� ��'K$Y�g�*�fK�\�%q3]8t��ז^H�#��a�q�##�?�X �NR.S��� `�9�3#lh'�vm���[�  5}U3�\��i���&"��1a5��F�`˹�5 XR/ W�����7�n � X!���
�iS��v���u��j���w�g��S:~����}u;y��N�R��̊G�-=����Crd���z���行���c����A91񈜜8��N�SS����19�q�f{zꨜ��t��'���:ǀ���#rj昜�~Z.�<+��:'������ݏ�c{�{�s�����Ď'�؎���N��{R�xA���3%���X����r�]������|��?����M������)�*����ɴ�ј�  @M��S�F>���oR��I��<������S��;LYk菡a�|s�.�%p��ѵEju���d��[Ȧ5��l���)�j(�����L�  '�0�Z��/��`7\�	 \�`)T0m�P�0�)�h����q���@H  	�uL�k�x>�cKUm�e��8�-Q	8TLSR_1-�@@0�V�U:\sfH`O�n�s� `���[>0�y������@��t毝�0w��;����y l��� ��z�ʚ �|�%t��ۺ�	�fy�tx�Kp���/����^�G6�� �*�[�M��$Hvtj�D1�^���!�xX��1�p.��1Y|����c��j1 �q�_, ,��1���^K$g����^k�>S�毦�5*=�[e�h��/�K M ��Fד�_˾k2�: 0��7�_����Ó���Y����<'�u�ߙG�����Y98yJ��O�#c��p@�>֑ :�ᱣi����k����I�C��8T(l��Y��I9:s��x���1��>>�t��I��!�EG��'��������:��1���3���ӻ�ltj�3r|�rt��rd�Wؾ 'w[S���M9}�w���?�s��Jξ���;�Wο�W���PJ;> o�S �&k0���I)��,) � �R^;.՞)qy����oZ�> �?%a�q�{14�?��:�-pPǾz ��� ���G6��-}n��kL-�����_�YP����L���혭���_t/[����Lq�^i=W�!Y`�h3�|-��5 K@�` ��� �P�%�:%���'И�+� @��d@��s���"\��˂ ���#�ZZ�*>Sɹ/���� L-@��� ]�;�˵Kzk�H�G����fh��~��!	������M�+�wc��*犭�3[�P���S3O�����>����Ok.����S�l��ܥ�Z�!5�[׊%�R��)�랾�����>q*e�� Ϻ҅�:� \�� �0��о�r@  V��&�T8�6����^��k=a��Ø�*��1�
�c��q��]��@&�Gj�-y=F͹��ۦo��5��0c��q�_�?��+ W6�ϡ� �  ��j t�u ��r�?�$oQ��jy&���-��n��v⻖�2��:���bi�?�7�_.���r��oW�� �Ko�<����?q#='G1�c
������������ɡ��r��y�|D�9$�f@ph��#;<!'�`� �6�wB���q�c�ϒ��~JN�fNˡ�j�G���I���� �?-�����d��v��c ���Sf��1���!�]!�Q9���sd��vrC�|=mt�خ3>)ǶY��xV�����Љ�n������r�ޟ����Z������;!'���2�\7�ny������!-q�K�kҨ��Ũ�p�H�gFj����ϊ׿U|�Y		,�Y��I�m,@&韖P�D
 ����:Ϙ4���m�{ԨA���eԠY?�_����t19�l���c����?�,>O��c�(�r PK�s|<"��.��tK���]mR �i��n-�c�>� BF܃2�@�0v�0��`�T� l˘7��R�/�P�i �@��J���Z���B�v� �=9P��騀��;kvH{՜��̙Z[
-U����5Un���Y�+�F�N)�W<"��!E�| "o���ٚ�	�"Ȼ	�n�����-Aֳ�E���5
r�u��`�t�`m���x�
�!����J��N���l���8t�A���>Lȟ\䫀�1R��:��^۰���,�h�G۸7I]���W�=�A6m�e�UZ-�[EW���!����������]�u�v��=��s��5�oP���(�'I^K���}�%��%Q�N�p�v4��I�5+A��*���s=}�F�4�����a�r{Z��GzO�=R(H����\�n	�b��ĳ���E�
R�Ta�k�G��*�d�`�ŝ [Q�4�P@� i?  ���g2�,�����t��ϛ~����l�0@���#n�ͽ�fV�p��2j�@���� /t�1 ʁ�u��"Ĥ�j�_U ��f�/ \�����J����c �9�T �'�?>y��M�����ә��N����Ԏ���~G~��/��B~���}�����	9=zJ���W��~y �:&O���|�C���I�ѿ�DN��7��}������L~��O����G~��/�g�ݟ����񘙍�	 ���8���;GO�������۟6�' ���8 p����~.O��+y�������}���|�\3�^�n�ykh' 0!Ů�% `� �Y�U ���6 ��4���9����$���iI�T��o��
$}Z;`54�F�5�&��#�{F2�wK P�4���  � �#5m j� ڌ1y0(�z��� �  ��P���6�
 �+ � # B @�@�T� �d�
V�K�\f ��@`C�B ��)�KC@Y�@�k���^@G�`k p���ũ>2�>L���ty�I�{���w��m�T�����P�o��o�R��x�̕)�m0�)��q�bde5wtl}���W��/My�1_Wb�(Mś�1��7I}�F������K��F��B�(Z��x�Ke����b�D�7r�7!}<Ⱦ!IVr�U�f�h����t��N��.��o���vbؚ�_�l�o+��;u9 P�����h��vv�߈ &��.��Sh��zď��1}���-�= ��t��0�NMV����?�0� 1e�5
 � ,�;Z `C��8����F����?m�)~_�?H&1�8���?D�P�/ ,������ K� �~�܀���{�J  �7����1�,z��t���]&ע끁^�� ���Qyxb1 <*ǳ蘙%��8�@������<!����W��5�P�z\�8𔁀��}\̊�c����|����	�����#��۟�o~�;rr���?��Q~���C3����'@��;��Q��8���'� ,��3�/�����ɴ�r ���Į��N	���r��oə{�/����<q?���ʧ��5���OVmz�\?���m�rsx����k� |d��J(<'>�Xx����$��$p�佩�V`�	_�B�����&���F �V=P��C�  �U���R�=���t��K ~��O�S]V��b�~]jy�}e��!�W��2P>&A��S!�:���_=��k*��{�(�sk>�y@�Y��x������iv�M:;���6�V�^���f�:�M�g/ƸG�\;����m�P�ѐґe#�Ώ�5�hv���<�CW��`�Q�_R9}RǾ�\̟� ��U�8�< R�:���Pn�h��H-�@ /�'�* �e�3� @�lYn-�l  �W h��_������=p޴�x���ٕ�b�w*��;�� � k	m���@��l�7b�*�����)3>ʎ'�˔!/��Sӷ���W��Y;?�ak�w�2� �
^�Ɯ�}hS�B�6t�Ό�����l2Ɵ~ܰVe���I~ߘ�J�e�Ĵ�)m���d�(��E�ċ� ���  ��V���:5o2x�C��Qc
T�ؖ���ƿ�U���oo�7�k�~�:^{p1D����q��<Y���Ӻ ��
��g��i a�:�i�@g03�٧!���UyPi�C��c�/�H�Ξ��s<w �J�
 ����#�����,�{h89~��?&��~�rn��S8,�Ǐ�Q�Bk����� � ��{)��id���=q �=�-9{�����,���r��ߓ��OI��������[F��.��LH�kL�1��ک�� � �.�� `��";   4'	 �,�Y 0E�B�}]`B�Cd�H���IiA !0&u�Q`aD��aI�0�����K$D�1 �"�,� ���|y�� 8e��򓩪��J�������[�]��0r�B��; @����<n�WPH�d���5�� �tT��0}� ��w�j��] l� ` �?/��Zee�  ���_��DF H�c�:Q�Ώ��̚���Q�S�,2��D0�ƯR H*   �����y �����e���ՉR� @�{&���" � �5 -5�z�Z�}�Q��4 ��w/�nϼz_�w�t�ԎZ��Vε :�OU�����-5[W
 ��3�a�%��j 6 ���w����OF��xsum����U Tj��5 Aʜ���1b�P �����T�Gu����N5P>UN�_J�{U�Κ����2��_�1-Ǹ����5 ��j�� ��������ӏ�g5 �U�VY���mp���V�#���T�;�-��'÷���L@��7���&��ްZ�ɂb�'&�:���y��19��	����}��Q@@����������g�RN`�f�`L���	����w>�]y�����Ͼ�9y�}�f� ����G�������[|�!����/�w��c ĩ1}��( |�rv�Y ���Q @']p\r@��n;o ���c�	�SH�_ub�B 8 � �����G�w�a��[֌�/�N�Gn����:�!yK�n���~Ř�B@1�S��kg��3+�ޭ ܁m�j  ��.��X) ��6I�#`��$��dpF��I�� T����CJx)LH]pX ���6�d�dt!�������W���@�& ������!�*AS�b�^LŇ�{���ٟ�/��ߖ й<�>�:A��H@X�*��� �1��2�幭� x��LW��b�Ø�5K�N'k&KR �x�aޯ $��%U� 0#Gt討��# @6�����& �fϔ��݌�o����ܻszL��%C�2d����k �;5U5:��F���]��VV>oжԸ��{�����	)�V!-��yuH�5 x�T�K 7�n��Ũ�W���rB3����?��)��i9�ЉYݧ �8f�8F�0��xR~����!2�Ó�J�i92zZ��Cd��}���}_Ǵ��s�~A�y�B 84qD��������~D����ʱݧ0�#f�a]s���a���~ gvi��a� tD��i��	�����s@�.2t=nt�}�����L N���<z�7��]ߓ����|���%�~���K֌�/k��++�~Dn��Q��u���O��v\J��K0�L�T��k��Yq��{�s�'��P� ��û%�-  !i� � ���$��R�Y�F����[��"a*1L%:��0��8����3&	�&�b��K�N�6�p����v�� Pb����U`���Gŋ�xj&.+7�S����PpM��vJj1��>Gm@P0� ��v.L�I �5j"Z��<�y�  �� � tN�G �.����,  ���o�<l/��n��m4�i�r�]�{�F;ޮ��iQ����-�
]�ӵZ=�@��^��`c�OPV�%�(�Ns_J)�V����.�[��+�k��j ����a�+��j��v����F:��<Fnw�˪��IK��h��ke�:h��i��f��������v���8-�}F�ݏ�O��Wr�=������a�ڛ��|��ߑw|�4<u�s��_3�*�xh�<������M�>"����ɩ��x���V|d����?�ӻ�	 h`�! �,H4�� '�  `挜�j�q]Bx���I����cF�8���m��_�㻀������_��}W.��-9�����]R2p���[�N�SVo}�,��Y�������.0%5�))#�/#�/�lM���%���?f�n vH �EwY���l�Q�����+��[ P0�G�ƀ�Ĭ�'y�RsF�u�������E��.4-u�ILM �K�����ՀD�0FO�w�S.
� T�@G(hg@]Ԟ�i�t�3��Lۿv�$�Z����c���*�:s�Hl�J��:�2R�wc��*�$�y#W�gj�=n�θ6 �d�ּ\#/�櫙2�@�&1f���z�4�Ghg�N] (�����[�?�= ���k��Oz� �V[�t�?ߋ��h���i�ב%@ f��c����*��D
6r��y ��$��& �ۋ��K�^�kN �!@�ի��d�Ɵ�( -�X�n{�6����En2kF$��Ư�4Et-��A@i��4b��n��Q{�8��׌t��b�
NwZLޱ�"���r�A��� �l�P#� �>#��֥  ��W ���e�Y:.�b@�h�A����^`�"i����)��
���:�̹�v��,ݍQ{1m� ��*P&C*����b<��A�L��/R�B ����y-���Zj���m@� &*5cK�x�����. �G��  |V�e���f�!m�O�ƫ n��� О���;�z��_'�n 2�)m����܏c�'�����l����A�ض'�0�����D����L�0&�+�N�{�ʏ����2�O�<o����Ә�Qyc�!�?��O���������}_N�8+���v@A���Q���PN�|��18�C�xM�� 0����@�q���	�q^ ���/����Χ���g��m/șߑ3����m��T��ɺ���3v���z�����u�Ge��ȍ ���4Y����髴ڿҽ�}�����3� �� `' ��� @� ���-�`�1�6 @�������@%� 55����X�C�v56��9�x�Y� ĶJC R�	I qװ�&��uy_��n��Z Q6㷵4 t�� �h�6e�'��M�P7@@{Gk���m�^�ě +�n��6���� P,ԒA P-&��Z�k�����ת���.���:y1��v�(Y=e���BA-�v���:3��Ew��Ig�6�	܎��.��~�B�����y?� ��V �ٵ�@�����)�u ��k?��߬�H����0;������	� 5�z��� ��G��񧥓��( �+B'�Ҫ];Bk �s��u_
��6+Zꊍ���I `Z:][����4�?T��&7a�j ��ԋ ��2 �	  @�s���/���c�:y��u�2�k�(KRx�
�K8��|"/�lA�6X `w
�b�*5c5����������� ��g��^4 \T�( �ʊ���!�|�1 ��y . ��f�Z����^�٤=��������� �?  �mrpf h毦���X5g��"��崞&����i�ѧ)�����O=v�W��S~z�W���o��ҿ��W���#y���ȓ�=-?��O����Q 8&�����85zapX;N�o�r�
 �� �pB��c�.ȑ�����'  mxJN�yF���������]'��*yݳ�jh���-9��[�|DV����- Ә?�?�� ��@���� ����d��0�&��d���5�W������ ,�Q� А�[`�͍��Z�wKs3����Ni�ג@ ���s@@�v"40*��a�TJ�`��Z �`j��i�R ���kL/�M�&  )xlY 4�wp�Z �ąyUb�
�wհ�	 �#��x��n����@��0�P(q	 0�� ��?� t ݨ�@���:Q�����̥`F����BG%��9�!v���duZd��L��� �p���� kv�>����a���F�^� ��+��9@� �� ��e3ע��LX5 ��N`g1 �$J����T. ���3k�L-c�ֵ�[j�t ���ܘ��Vqc��K��*��[$yr�y�׳���� �� ���o ��on���V����۽�u��e����f��n����_k �m'�~BNn%֞����a��/��s���g-͡m��ѹ����'�w��|��?��|����;�)/����د��"�� ���rx�	9wד�~�������،����1����;g�`����#�3N����w���fD:�БE `�@��� pdۣrh�crl��������e9~���w�'��-9u㲼wFVn�#9�wʺ�������;>(+v|Hnj�f��J�L�� \��f�>�F��[����G&�Dt��i�`�Ā5�(��
 �	0��� ��k�o�����L�k�+ͭ� ��<�+-�{��H�&@�A��3�Ԧ ߸�jG$R=$�
��x@<����hPZ� `��bFNX�\��<k� ��Øt���  � XI��u�d/f� '8@���rk��H � 7����[M���V���Z�ɹ�������f��e @�G��ͷ���1|�����F��s@�����=����i��!mUs�Z9k��.��14"	LU��u�]� @��V�N$�<Z �1 �\�0`����s�� m:����$ d���ִ�����TH+ �ʍ�R]�qX�8f]�������Uc������y�w�\P�o��F�@������Z��6Ԃ� f�Ј���-ՙ�_: P��`���1�b��B�5X<j�����s�@&�W��1�o���I���r���	 <v� P�E�ƮR�u� �1�Ĳ��f�/V�ep�^y � ���g�u� �  mj���%j �dӛe�v���  0��&���s  F��ߡ����}Nۮ��6��e9J6}d������r�8��1yx�99��Y �i��Q ����[����S��:)c揨0v3���1y�P� P- ێr|�crr;��	9��)y�Χds�]���ͣ��{F�억C����e��{�����s��ȼ�|S����?e�����\�i2�  �A
 d0�0�Ѭ_'���� �~� l�W�a�m����҂Z[P3���z2" �A��3�C	u>��gT"5��Ԫ���)$K��k0r�h2�,p) �� ��_o�E�G�8i�� ���� ���� ��	 �Iq1���7�Z ��� η��  d�Q9�% �����{e"x�̄�.[#�m�w˶�{d.�^���dgJ�������\�=�5����'ӑ{e<t��o�!�m�����o�8�����1Ip�t�D�(F� �|�@j���� ��oC�1�E ]� ��� @	�x$Kt)۴��&�������t���fƿ& ��|L�QK��I�3rڐ�)ѡl�~��R ���J� / ���l:�-�� �Y?�k���� ���1�� 8�K���� �eԥ { ��M���> 7�a �: `�Sf~��;_�c���@�阾'��ہ�� ��{^N�v( �>�������y�\��a�lUG�> <&��^�C���I84}FM� ��1 `������q  ������3g�ً�>6����8N�{9�;��{F>#�Um�,�#�4��)Y߳KV�&�G�e��_��> ok�)�^L�5!�	����jd B�j`�)���%���@��^��I�o)�E0��g�D�3�x��� �������n���ۥ��viEm�mf_�>i��i:
�ŶJ*<-��AoL"�	U��l�x�7H-�P����k�$T/ l2} ����)����� ���ymP;hΉ�s��\눀( g�t�N���+w�}X�c������I���)�,���i����������Y�*ݧ�9.�;*�="�F�9"�1tH>9�0zP�}���o����|\���$�� ��+ �5�_� �Z*��@�汎� P�kt�zr�s��Ë���n1�"�d��-���d��$�G$�g)�?�@œ/� ��*�_Ej�y�{�4�O ���k�(� `��y� ^f)���6I�Ƭ����h14� ��  �}�_��+ Y p�����d��Z�& ��x�Jy���� ���O�!���G�]Ȍ���_��1�]i�~���:�2��c�_�c�OnVNl����}Ft��ѝ�.W��g���s���횉?ftd���vA�����n=%g�:��198q�?$_�<(_�>H`}X�8�0����zD�>���3��)0���C��j��C�}x�qyd�q9�p�}R�R�;��o��Mrs�Sn��(�[�em�6Y6�G��!�F��%+��#76n7钿��S�T�ՠZ�Ů��=� T!� ` ���������	c��1�%� � ��h�� 4�oo�/��I+ `�[��v�@@�m��!u|6�*��$�1�o�J�zD��[ ��RK�w���K�)�K� ��d ��oz�M��5 f�+ ��x��	 5�'@��k�rs��Z�?e ���o�;��<W�.��v >�AМ� ��p� �l �  t(ۮ����gN �@��i9<z@=��s���9��$��0�N���ZOr�?*�|F��J��>8rR�4<�/l9"��rH�0���gG�}Z��o1� �[3��lF� R9��;�{ 0�0�d�I��^߃�c� ��0~����F�ԍɣ�22�J�|]�n������|T���eK���
�e0v@���K6��|�T�XF
 
��/�)�� S�! ���`) q��\�  �7 0����W>���} �  � < ��s� �j��ߥ[���si� S`�� P� X�/�b�n�W �;rK�Dӊ9����i�W �Q �T�O+����C `A �2 ���M ��o���z���W
��u�ڿ^�U��|[o��[�MF����F׽�V�����m��F*nJCဴJ[��t`u��6A���+����> ݡғ�>�ݖ�~�
�Ψ3������!�dZY�Um�V��4�f��F�a����q�ߨ��Ik�i-�(-��D�jD���:�e���K[^������u�5�����F�n��.�+���Nid����RXT/+
㲢�YV��eu h����oV�m�#�[Cwɺ���uӒ�&��x�1�1!2Q�P͘tLK3W ` �,���4�g���B�-{_D��MJB;���J�Ҙ��f�z d�m�a����(h�/�ͻ��a�ԥ�$���DdJ��q	a�!����oW���h�B��z�zm�T��j�@�2j Rk��@�	��N�}�� P��  ��[�ٚ�c�Ur,U���򼘰-��[`��q�3Rժ�cN5cRU=
|�I5纆�V㛒�x�	o�_��ׄvf�
�,�{f9'�X�$��Sܓ�ۤٽ]�4��dt�]m#�?��>���g���yc���?q�W����90z }L������O�|O�� O��k��}G�0r\� |~�8:*�<�������𗤣tc֡�:�m�d�@UH��b�@�
����mP%�WS�:D <]p&�6�o�~��G��]�ޚrX3����Y�N�"R�����y������+0#�? �S�!rZZk&���A��Zt8e!��E5 ���/�/���  �ݙQ«+ Z�[[� �5����0��Y�ǭF��i�-�w`Y:&�ţ�*7�-����$����&o��Vq���V� ���P�Z;�Z@����l���	Ѓ�_	 �om��m�f�ތY�x����i�N�_��`^vGEK��Ok��;uy xt x� ^u� _	 ���ɿ�������/�����7d�uaY�֘,�9%�om��˛e97܊m�|e��X�)+ٮB��W���b�Z�E��|�~O��i�ϗ5Ȳ[�Q���o�|S%�cr�["r���z���Z���&�����r�?Wɭ�T!��o�,��RY�Kdտ���-�UoDo*��o*1Zu���3ZsC��}s��Ck���Wr��| (gYDV���s��>�Y�;$��W�k$߳E
#�����6�i�.k:w�M�1�qKm%�C��Ѫhɣ�ڑ��1��{R��S��;�?(ز `� @ԇ	tb�i��a}d�?��v�km� � ���K2�M|Oԯ��ܾ
2��EvWC�r�V�:�ڗ |:�@���0�!����S`��� �9o�/ ���qL��)���� ���_��~�g�~,��>!�������<4C�?yL�8yT������? ��
m��}3����{ͤAwO~� ��&���wI_`�4q-�d�Z�R��5 �kD�G� &���$Q��Zp���lf�Mt �H �{�� �f��onͪ�=�m��on� �  ��+��)"(��Y�#�X�x)>�_4��3RW�աIMgTW�I�*7J��*�T|��E�-�J�ߍQ�BE�f}m�f3�\��<��S�P���6���y�;�]�*��6�aFț���O�˨�G�%R�d�CQ�m����w�H�5��}���|��$b�[�����-9�1Y���-�(&4bT[N`@��Qc���a��Ae��#Ȍc�F�bX!����43�z�C0�s�S�#�@SAO�0���}Ҫ� K�^ `7 � � f �tmٶOa�x���� @�h��6 P���! �O���� 0��#�����!�Z�ޒ_�Q�LP�r�iX
 v�}��&'/�������<u�W��m_�����<w�w����|��~.M��/� ����������  *}������f�q�kx��'d��^n�]Z�F��-2�x�l�z��s�săqI�[��/ t�v�c�N hD�g[ϵ���^�����w��Tc�Z��_ a��5JDuS#АUN p*��۲��O���}��u�^+oy�[�M�{�E p�_c�Y�&  ���ֵw�\��[����B��s��	�ڹ'�?D�� 7x�=X6!��I	�͈�|�l���MK��+�n�
�����O�r��o�J0�BT��G$�;H�r6�Y3�B�]�'>2T?*H�
�G�B���_|.wAm��7��K��
nȈ)TGa�+z8�-Z3-	L �&k��@d޽��q2�]���dum�Um��	e�	DF[��ܥ��Ͼ@��* �*����7
X3������;��6�T����΀�:	���5����m�-�:,p�44�:�%��)��v��`s�r}0S/��<���ѶK��� �[�g���| l) ��.���y� oa?`�[�JW � ����2w�D����6����p�jj'��;i����� �����*!� �T;��l��EM���˗�C��i��3��yd��8����w� �w=!�&��w?�3�y�����<2sV����|��?�/��/��4��� >��s� Ω@]��/�l ���F�毊��Rz��- H�,����o! �ڻ�CRǽ+�d�4��8A⠝���?.��8 `w�;�V`��/���+-' ���KjF���%��$e�R ���� o� 7��C�R p� �- �� ��[6X0 Ls�k�QZ�V�Mk� �Z�T ��f� f���1}�c' �����	 K�\J�[�}TK �-]�8��f��ty �  | Й ��U��U�䳯�N�K�-r�_-˪7�Z n���Q��`�bPby���l=T�	�b�Ә�V��Yo�j���l
�@�~������� �o֖LA�P6�MAsSм���f�@��%��_��$�~�ErJ��e@��8q�q  ��&(�I�'�ꀏ��q����Y�\3��:7fJ��JAU��*o���>qo���M�M3@@���c]�FkU�@� ��H%�i�	��BU�s�,P �r��a{:�O24%�ȴ��Gbִ��7�wIS�in�k����Uuu��.I�vH<2'1�H��+��+�L�&=���A� ���^, ��y� �w�Wh�	��t55o�0�ނ �Zl�/ 8� �-&�?i�� �����F�994�:/�xA��='_}����]/x��(�� C |h�礵�k� $L��'�j�d�j��I�l�x-��{�P �l���T���l�_�m������5�+픕m����N�O#��� �^�ݨMͿf.=�Ҝ4��ձ?��� ��djԴY�2u�&� �4I�6ts�U�Sٌߖ@^��Q�  \ ���Y!7�Ŧ}6H�,�`ᤄ�&$R2`���g��Y	_�"|.��UѲٌ"(D 00�2���~{���L��O�0Ĝ	��c���$޵� ���� Ѵ5�x��o�)T1U��3\��c�H���Z2,���S.���cR϶c�'㬫�!��J�@ ����ᛖܒYQP'Ņ��&X�
7�U�O��&��ߚ���.�H9��[!�gT���*T��<�c�/@<�D�%�j:��ꀀz�����o��e�k�*�$va��%�&Q�螔�V��c�
 ��  ��@ �ë�S1��`p��A񖌈�s��d����w@�e ��% m���)���aӳ� xx�?-'��1���_�v����NX����0������g��Gx��|v�����҄�, Id2Ԑ������`�Nk��8���@�.nP�T�˺Dq�h�� U�}�B�Cx�5��@v��_* h��3jU��ڠFTϾ:�b
�s ��� ���n�z X�?���^�WJ ��n��������Y�E����2�7��oo�Eo|�-��q���/e�怄Ȑ�d���		Mb�S��B����g�W$���1�
5{뱭`Z�����"L��䍡Q�C�z� P���� A�˿^��Y΂ �Ŕ�E�5~�z������ �8�co �J��l��l�3pYJԐu�d;9��e�������_]�c#0ۏ}< BV3�;��Y�ʶH�\���(T�P��c�Z�Z��3&1߸$���3_2�hM@���$��3���d���&)0Ծ:�k�ٿV�k@#��b5 @M���&3���`�3��ꔥ�0x
�[� * ��Ny׵qm�ş�ii=��5�@�� o�#]��sF���s=u!dU)����a������ש� ��r<��՘�kB���*�Tf�*4+��9���IUd�T�w��R�%5�]����gN|�mBQm� �h1 �~ �]2�K�����޾���� ASm��||���(���A��Mɿm~D>��a�ئ�c�������䁁O��6�������]=��w}D��������̑Q�U�i�I�t.��z��s�c��4���M�_M�_-��-@@K�Fi�>o,�Z�R�}���1�ҡ~��n���M?��>I� l����^c�����Qx�ut��X1eH@A�x�ڵ! `㟟 �7$)���E��\:)��k'�݅aw�v�Eջ2��.��c�-|Vk  ��:ʥB���Cq�a̳M��9��9�+ &|��b@@ �( ��:��ʺ�fF�ө��o���< l�� *b�1}���XTKL���w��6ҕ ��vJ5奆rc���V�X2 \�!�� �f��1� 2�i��B@�	b��
�8/
�Z6\J:߀*��]�$!\�V!i9��/�����@��L�E��T���xI�,l X��_�} ^^ X ��Nva  d@�< �K�%l  ej�B|�6x��/����R � ( 
�ş?F��YM  ���?����c�v@�`�!5~&(��j�:��*�A�T�q��8 �K��b,�6IA�Q��d�	
�@`+Y�s�ϙ�9kR�bM@���1��_��ٗ���1���>���+]*� �2@�@��
Ul�(R5$�j, �E&$ L� �#�Ŷ�O!�&�ǿ�cfd�:�P��yv[ `z�c�&�9 ��~1 �b%��e� ��m	 HC �fi�5I
�C��iTU:������T|�C�-6�:�{M�Mn���  ��j1 T* �g��W� ���� �m���@��Z�^�np�M5��P�t�&[j-�M5{es�>��{6T�����W��*�|�W�M�Ȃ�˧��t\�o��ܓŃh���/�}H��iѕ �d���f�]X��{� hr[��@���)@ �}� ���Ў� @i�ԕYj P+���jX���Q�kD��(�P�u �&��rB��'M�Y}�4�M���j4%md��dҖ��b��2ۗ ��U�  �_ �< 
 6�즧��>��r��P����I�j�a�k; ��<٦�T6 0� ���
 �����E5 K  ��� Y: ^Z~ `�֔�'��(hM��c�lA�$@�\�qcVa�m�j����jj���2]�l�'C!�L����vLR���\�5 N%P]A�\�*&�Vz�<�E�k�1�.L�������a���#dPQ�?ZA6W��Z�%�B����B@ŠD	�
c��	�z`%8-�ǧf�*�(�[�����S����v�����d�35U�_Q���le��r^_ ���li��i�c]C]�ؚ���)7�X��_8$T˾Z���3�% �/�l�������K/ ��� z�{�׽�>�m���o��������.�^�D�hh��%-.m��;�V	cQȌr"�7���J��T`垱��7q�s�r~yɪ�>�Gͨ�{��m�����[�қ�� ��:�@k� ���kz�^��*���~i���5��]�9���U �q/�u�@����^J���F�\6�V����<��)CU
[�d X;kd�@���� �4, �b����Y6U��;�j�b �\i�B��? l�R p�R`��k �rk) 0F~�U*; � x�?�������4� ���p	f| ����2����RZ �7! ��i  0b � �5 6 ���� ��-� Kc�$`eS�@�P�9��_�e+\R����O���XU!�dW:fZ�X�k�)�+�X*9�@-t58L \
 �C:T���\"R9,Q�7`T��q��N�kM�F� +A���<��__�z��d����gͰ=j��[�L� �Flf/s ��l���~����_u� � <��ER �z1=m��[g\+ҩW�,("�r���s��p @% P៖
΃�Yd �S*C��
�
����%@G$	�uu�����]ۥ����ѵ�1�N5�٫z�x��w���ni��Z1�V�����r��Y�)@��-�������Z������v��a�E8�� ��1h^k� �v����v�6����F!�	 	�G5|즀n�ڿ����� �RW�+��+ Q�o�z�F̞߮܄᫬%�S���aI*LsMR�@���&���|\Z)3m�h;e�,�y�j�_ :�wfd�����.�� ��Z�ӊr��:x ��� vS�B�׮�-�-t(��O� `�Sj(3*�WK9ʔ1���	 ��-F�� �U�c����n�� r���.�l ���5- r��b � �B��� ������H������G0�A	�lA"���T�;j g�V��K����ZҪ#�4���� �H���9+C�lY��������% ه(�&�j�*Y\������[6 ���'��W���д� @ ��(Ƿ ��(T� 0(a�%��G*1��1�)�b$:d�3!Iߖ�S�j'��Ca����>�f�Z�s�{ +5��@�  �+ /�i��pN�>�tu��Ц � P|�C+ <��p�_t�� �՘Yd �; {�> `�k l �\���62�N�f�Szjw[F�&� z����v�%��� �f�1���9����:��|BK'�՗p� �Ei��޳�6� �=����	�IL&��4`�@{�&��>��~��Q hMC@�}=��i��( ��j4�[�� ��Ti�ԗ�q�o����@R�@�����{ʹ�ˁ~C�L�I�����I�K]�6g c�R6i���( 4�FԀ����@ܿ�m ���{���E �] ,��M �t�R~�Z��\,R���R P� ��y� ���� �e�k   ̘�s@�S�`�2`��S�^˚%�3~� ��oe��z棘����z��VV�7"h��%���A � HI`M��)�6 �W���Ob�)�?��'�7�0��A����ZҶUͪb�J3B�,,�]�@G4 �1 HGt�d�f�@50��0��`Չ�j����J @;�i';�� �1=�9�^@J��� �'�Y��C�l�!� ������ >`�	 �!PG\ v: �2����+ ]���i�#��MV��ڃ0��}f�C��T7���q�j\m|�x�9�9fm/O I�$��y�z��j׼_�vCQ H  �|Ku\�������۸~�a'�x'��Y>(����  &� �M ��� @�� /RuqL�����M�I  Y�g�(�.C�(�)�c�q�:b �1�o�z`@�����P h��ڠz���z H���A��	 �lp�x)��ȬSܔeȻ�b��B�5�e@p� ��o���5 �s� p�_�ܒU٫��5�R��_������7�*�� ���X�ǽTP��[ Y��ba��u6�x-�{��Ufh &o�k�n3� Q�!\2)�2עq��c�]�N4�Ȅ)x
d�uXR�4C�@���%�U�f;h&3Q HV�U�9�n�)��;D���Ò{�_V�T&UkR�N �]� @�����	�I�H5u5w�nZ��FШ4�zL[UW�1�z�rH|H� X�����󿵹CsʹzX�/F��W�H�
 ��x5[L?������CTppntx��s�'��9 ���O�u��j�� Z�KA�)����?���@ @�[� � '�wM?O5`�15�����|\k���#���bT:&>�i��,d ` ���3 ���������n� *B{�3����N�M�W�=_��& � �Q��7�l3C�4�W �~ ݮ]ғ�2�.7����x t��v���g��5 ���S�?�S�l��ڐ-koz�\��v^�Q �$��N�b����\�F��f̶U�����Ž��=�U1D���A� 5�X5 I���L�ϵQX���� @�� ��@+JT � �K���KUxs�G\8�X���<�XǽY_4$�%#�\6f5P~�� �/�v�V�Ȩc	-UP �
���S\��PA�;�vJR
�A:�@�g�y8���^�x�KhЭ
fD@�5��}�  �HM���E"���-�B@-��(�������qp��j��/��DY�Q��fQ��� F����2��  �컥A|��/�� ���d���Q �n�C�F����#ie��U�,��c@V X�V�/�@����. �C��E� .�yT>���0@  � љ y�����&;�_,5}]����� �� ��+� �|v�@
Y* Ҋ NEK1z#h㏕Ρr/�y1�)�(�?����QF�� �ڜQ��- sF�Bk���Ɵ l� ��8K!�� m��o�� �� ��aɿ�'��Z*5 ap
z<�,	 H�5�����M��iu:�f��&Ԩ ���� ӱ
�VȈk- �]��i "�@��^�p���A]30�cO�a�����W��	!�ih-B�`��b�`t�Em��i5�1h��* Knm�|�-���r �V4Zp��7�@� С�*3ǃ���H;~j��?X���  �Of�#�֙*�\3/�ҽ  �J�@h��B@yx�wIip�T�k�N � �Z�5{.  F���aBۍl0 P��6���5 �yM����B��D�ۨ��� $��V��WL� �Lu̿���2Z�5`�M�kj�}��^�������Z y ��o��Gk����� �&�����i�$0�d�V�o��Z42��tH�� ҵn� ` ���� ����^5	 Lc�֐�N=�i��y�� i H  )L<��� 1}U`WF1�N#5~[W � ��� j ��-�����y]iq��S�)�������<yd���3`��.��B@ ,o1� �� �`�^ ,�X$?�o+  o
� P�� �. �倝Z *��N 8��<v��/  ɲ���  �'� h����� �] ����	2;�.�ni(�+���t�4�&��%��i�Ԙ������� ���1���1�dV- �/�&� � �]M!�Ȃk��?]�_�m]�F�+��oJ��Ϳ�l��vB�k�4���F�U@������Bk0��θ �>�i�����@����[�M
�®Q0���^{�6�s0a�G��]K�J�`�� S����K@  �J�pL� ����@�����[3!.�k�gZ*}[1�Y)�IEpN*�;�����	���B6  ״�j��pO5�ԌQ�a>���mH� �pu Pg����=+�M�f�&��&-��g�V�u;��6��q�X�O7�QG吴�oY ��z�v�+��"�S$��{�������f��=��Ήii3EX���7��R �P1C9����HJ��\% $B{$��ٷ^ ��֙/�u��Q��,_��u���Q�
[x�[����� is��0#  ��� x 0p��j��	 N�����k �r�O ���d:�e���� ��d�� @�IT�"P씞�����л��;���lgNR���q�T �w4 �k礋�����  s��^� ��z5�� �@�  � � @`M���� �m��d��d�:���ϴ  ��}[ T�F ) h-A#p���Ǭ�o�G	.jj����@��'#L`�	L��w <�*�!�>S��}
���z�Lsߡ��Դ��B�o5F��m^�N" (B�ܧd�A���k���i-@�{Z�<3*�ۤ� vHU`�T��k�_u� �ƒ�ʅ ��@��% sm0U�IDky�^ ��ݑ�+ �r��b�
 ��Z�+���	 1J V�h�o2~� K����ۺ ��_ ���@f��%  L7, �� ��U��E��Q���)ź���t �R	�^L�*B��/�!�	��  � h�@� � < �{Y��om7��ƴ=�K)����P X ����+ ���q� �+ 	��C�R�[�o��R���SQ�����VLj�(Q�CR;����н��/��������W���������xJ����B ���>�h���V��� ��
�ԧ=��2�&
z�>N˼'�f���l�c�������2����˘�V��Xk' 4�����/ j�� `�Z��&=��LbHR%���N	�:�1�(Yzd��V�':���7S��$E旴��2U��uN�1BvX�w0C�9�4~
��A"Фu) 0A�H;"���$`.������^��O������  ����\� ���y�.הT�*ϬQ�w�@;�.�^ ��G�b�����	P XZЉ�k�5'�c�g�������Ͻ���(35U�B��TU�q=ͨ�߆��% ��?�W������V�F�w
��G\�Z���u]��� %;� Z�oq�q,��MK��l�کK @S)�>��bj �\۲�	��N�
 �r��l��� fU@�n�� @�a�/5 �r�t*p������W|�G�n��.bd7�-eͨ�%d��b2�"�R�O�� ��V�EzFNʥ��Yތ�7I- P �n��ڛ�w����ٕ��U>t�	vSA薆
����� @~ �V6pJ!��|�|䶏ʣ��sg �� �l+� Y̼� ��	��BEy�R PW�K�c��/��|z�q����>%?;�?�]�� 0�`oM3@� *g ��S������mo�J���lh��
 u��[����rL�B��]- ����h-A3F� � uڇ�`�+�%��<̟��M� @�v8L+��J �)Q�%�!��$�5�j�LV�'
 A  ��@��P��l  �ƥ�zR�k��ʀ�V��j�5��R�ށvf� ��� ��M�P3K�ƪ���U`C�0 (�`�
 j�� �wm�9��^A h���FΣ� �a�I�g��O t]��W�'�Ժ��  �%�1�?T��W9翼]�e!� Ŕ%mH7x���Z �2g&�<���e ��5 � \�٤`���U������� �  @�1���$�b�� (Ѭ��j���o�
b� �e���%��*Zj�,�$ P_�[��_?�;���S2P�O�}����i���ۯ ��  �3`RMU���1�#����K@��̰����+Ŀ�B��� �s��+u�2�F��sj�7�*G��mc�����Ǩ�z 75 N �aU
 :\R��]�/���luMxkZX�:ܫ�t3rШ�r4@`������Ȫ�Eal�@��Bezc���#� X ��  /h  � �j�P���,�P�< � �q���:��b\ܕ�@`@`Z�]3�>@0�q�ڳC\�Z� B|.��uJh5��J����B�>�Qi-� ��Y + �qO�� �2����rj�� � X} �p  ��s/t��
 ���1��
�o�8U
��A `�� p)s�\�v��Nd��r h���+��1�zTǹL��dJz�&%�I'��po���� � ��"@��y ���Nɵ�%�d �����/��K{1�	�wK��G"�l� /�v ��(Xf���0�ʛ6�f�
 ͘v ���������_ � ���&�Ǧp� �Q� | xRΟyB�8�ek����U h��9OĢ �*�k �  oƼo � ���MY��  �꾫��N8-]]0�t�A՘�v
�N�k�lK= ���o���Ig��#��"���%�O����*�C ���� ���M�@
�J�^�ԥul��jF��M�<�\�KIxYL�-a)��%���&�F�QL4��k��<�����T<�����gφ֡���T����iJ�A�'[�+�Ն	��ߕ�%�_Op��@@r}������:�f[��U�Ќ!4cM��̠���(�;�ZS�5�oA�E!F�2�a�k�B���ou3��d���^��iM��)���"'h�BK:���d蔾���udM��%�^Wz�̽�����M i)�P#�	H7�t� �,��jҵ5{�[A`�[�۳U<y/Y���`��D�b(�I�a��q6a:j�֪Y#��Q�� �#�fK����Zͫl ����y ��j� 謖��s���.�[����Myװ�t�tt=��� ��׎�E�)�A�s���ݢ����9-��f�q&��1uR^�N��@ ��1�@�f3lT����[xͪ�� �NଁdA�h'[WuP���g �Y ��w��22@�  p���~���I �R��s	X$��F\�d�4�?+	�vI�wH2 �wK%"�%e�؝�]8H��z�E�/B��p���;?� 0(�$��X׮�� �j�����{ S5~�e�m����c՝E��.��h�}�*��J즀6��#�#3���^,G��6I�ٿ��)�U~^�Lߖ��o���!]~XW#tʬ�Vx9�a%@�E:���N�k ��&i����\8�,zJ�:�$�����/k������f! ��W�T�K�u� ��<�[���!�*�K�3vP~w�� �%3I�	A`8��`��ٔ �P0�0!������7H=�ԔG�U���a�|���{�+�d���VMK��A����A�D����uC��Rd�udũ� �Z�l 6�@�E���D;}i��a�%�.mr��Ԃ)� �PG��M�1L�-.���:���A@!�� f�gZf$HZv�����@2���5�4h� Ur!7٢���̈�� \�T��q�k�V��T
��vS� �� d��\L'����̱��I�m�m ���gV��  � �dpٿ�L�@��6��w�n�_�sBk��_͟���k-<�  t
`�`����?��;��d�(ZՃ�wK��s�V����Z�]+��<�0��/ Z���;>L��4zL�8��\`{����ŏ~I���j���5 H+��;�R �V��ϯT�`@ ��� `��C�ۧ~';RHW�]����w��L��[ ���Bи=*�`�_��鴥�bL����0�p��b&�e@`1 h �Z�)aL��� 6I#�אO .�|�0�qi%��L �ѐΌ֊Ѵ ���VW�k(5˨���\ `u- �f adc�Fi!�  � @��V�nn����7#S���Ф�u�8 @���&@ 9�B��>
� 0H  �u�a��eC@�9t� 72����6	�0vi� ���G�x�r@�k���Zݬ�cC��� 0�`A�� �H �=�u8�a< @� @M#�?`df�d_HG/d ��! ������ �� �͟s�$ � ���B rM  � �6W�� ����~���Q�;�����5�p/( 茓*���  Ƹ(���� �>�W�sg����Õ\C�?��E1�X P�9N+� j�%R�X ��R�e �ͩ���@�<p����'������� ��'��d1�դ����!M / �l���� \�0@��/���ҥ ���W�"K�';Z?*�}���-�>i/�S����I���H������B��Ȇ l�P�B� K����� �S��d0 �]^k0��Q){[@��Z#����Ϙ�v�3���6��oƠ� �d�d�dA��f�kKᤴrnۊ1�C�A�[���V5��'�����`L08���� �j���MR�f�4�;͹>��t 6�̿C͟`� `KA�@�NJT��@��8!@k � moS�w���d�U��ˢ��̿O9����e  �yQi�@i� o��xD�d��V���@@���6 ��Z �C�gg�:�k  �z�bR�*��Ϙ�$m��k �@ۨm �a@e�\��k���(�E 1P�#�ܾ+���Q�A]@��p� �N2�'��c��1�� `�c 4��� U��7���NlO��������,�m���m�<�q>j! 8!���h�P����DJf2%�[ Q���X �  ��I��.�) ��'��Nb�mFQ/Y?��R����@�dTj�� ��^�����M����9_�R�I9q��/�`c�1W��%	wGF��v�c�5-�F� ���B�?�ci X�$�,� ܺŸ��i��[�2���l `��7e���;u) е���N�k�hB�$0�r�ȝr�ȓ���'���c�����?����
�n�Oix .�� �ѳ/��U�K�RM ) ��� ��^��߃A�)wm����I���|�E ����E�A�AX�,Қ��r�0"�4��H�~ ���H!���<����Kb-���S�^G�~�L}L�8��y�Ғ?!� @ᔁ�V·��sҌ����"~'c���!�_���$��  �Ƶ����Ж?(�L' ��tU�a ��]3!]���TК��avM��`�����|vf `As�v����W �&����������ǽ����|25�5\;#�t���*  ����,�R �T�iP�R�r��� 2�{!2^��w6���	 �aU��֚,]�p֚/S��y\ T �Cv� �1�Kq C� 2�yv	�6�H]�6�KC���L_�X�?k�n5�xf0������ٿU�?v� �Q�3�HE�D� ���`� @��?���(�n���s� P�V�^f P�Ϧ �-��-���ϛ�S��_�b ���_&�3�k��r��;����=����;e,L\,$�s���L	��Ix .�?+ h����y��ػ���90�i���E���M W
 N-�TNPpjq?�zN}鰔��'Eo��*
�\�@�kȘVm��*.�z
ӮǼ�K# Д3J��VV�@簙�ۄQC! ����3j��Ճ�Z�ER+���~�� ` ������`LzȄz�'0D&�T�Y=&m�E `C��!���Y�0���kٮ�0�c @ Hp�T ����9�@+�~Hȷn�x�o7���Қ wɘ%� m�M��Х^������R P��T�ၯ& H���[��A���E� ��]���{�E ��S��s���?U�r/G�� JTOb����\��& 陓�{�����g0~b
������3��G� |�t�s.�*�3�p����8�.��3#��Dm���x�� � ��� ����?�o,0��	 ����w�d|N&b32���ȴ�Ƿ�DhF�
�7k }�� &�z��}���W�������J6,�7 ���
���Maiu*�!� �)�1����b�S�h^Q��X	������}�$�椾l�4��}���������E�A��]�����3<�+IL3��E1�0Ơ�U�j��ၶ�M��Z�H+J�+�x!&S0B�G�[��@SG&��-�v�[�RpC�xVQ�0��j�rM7 �+��dN�7HbՀ�V�����}X��K�Z `= ����3.�y�|  5�Ր�r'������|~�� ���/�(�+7K�-Ҏ�u� }�m��
p�I�{Me� t׌cc��@�	h�A9PO�Jb0j4�@f}�D0UxFO��.� �� �����̨a������7dV=3��uhZ/����U�ڈ	n�z~\�\K�8�6
 E�A�*�R�:lP�׶�MRKP�-�Z I;* h߀��T��ۘ%f�6�X9F�a%1K�͹��tS@�J�* N�cכ�u�e�����@�t�Č�&I��{0���M҆)�
�=�[����G����U�=Q�m��g)�`�&I :T���_� ��P�_#ˊu �Y�l6�m	q��^����<�M��<G�(Hc�u���ٹ�n����VΟ6})�U P��[6 h%^h�X�6�q-ئ��	��OI�Y��!�:���εUR���6 �R�=+q7�?�vZB( 4�� ����}���|L<��Yz��-2��1[����|%$S��b #߀�1u@�����N�������9&U�$ݘ����D�1��3$�LT�S��;�]j׷�k-�8]+�Ņɺt.   #L�R��ܚ2r�b�~쾵N<�g��
�
��B�������*z��ח�hf�2 `�^v_�n�ж��L��LhV��68+�<�
o�Ƽn	�jJ7I�d��Wq'@' \�yg3�Kii �Y�S ��

0&��h���  � � �����-��3� �o�7�DF"�KG����� �x ���_:��K�o^j�K�S:�pT!��چ�yC1F�"*|�Gr�-��:���F$3"�@t�
X�A�uj�ԭ"("�FL]!�  F��ҭ�I�?w�'��S  8 K�2�-i X�I���v2��EG!ƎI�TLHw5 � ��~�tF}�S��u �����i�(�81�l��g�� ,e3�_��� Й� �9��s  D  �݉x1�e<d���\��l P��
 5d�&@���j ǔj� ����A?
 A3UK�Y��dx^�y�Z  ���@6x)@��kT��4([1�������[T���N�p�k۔ |o � ��X  ���4 l"��/ �!�S~0�[�?�t��6�-^
�b���se�4 �O ���P��R��hA  ��7��)�S5� �<�$AF.b��`�5�R Ѕ���� ����( hM��x  ؀qk���?@]M"Pӏ��9 � �H@�" h^ � ��V�Y `���-R�����l�:��dT�eU-�o˽�>#]Yp! X��b ��+�. �9�,ވ��/�B� :�p �^�%�G ���b�wjI ���*2�� w@����ȳ"�� @0���SM�RR P) �`K! Y�� ��z��\Sb @k �DM-�*Lse�DW+�%�Q[@��aׯ F� h ���&�1w<�:5���  ��e��ߺI�o�&��m�t�   �P�M �.���e�3�Q? �皔���	�N�v-�@ALg�S�(�� po:��G� � r7�.�j���aLN��B�� �f��j���ڪ��<�Z���0�L� ��f���i�6KO�tWKW����j��+  �4 D1G�sC@G�謙͜��m+�c��� �آ�c��0�BK	�\ϥ^�4kb���
酂l�7��#�Sfҧ�f�j������� �z���v��*�� ���L��LkuB � d&�`Y��k	 Ѕ��d��˚��(������J_{ �VK����ߖ��/�K�?,�  � ��_��mS�֫�V���������� �@�'M���=�^r@n����s���i�
�L�)5{���)�l� gm@�(]+P�E�sɺ7�kEJ|�� Z0 }_N�b#�	 ؄�o�����?@}Θ4�� ���d��C  �hX� ��5  0��9��zȶz+&��`�����h�vZ6�� ^�FN ���`�|  �����	8N]) ��P�� ߚc��,��q�� "w4o��G�k��=N���J�qٵz]� P�i�bVn��s2�K  �	�j�(����Z��� b �L���^��	CoFM�����Ι ���� ͜���b@�G}? ���mA����a�|� � �U� ���!k  Юs@T �z]K P���`�5�5pq�y ���RF14  �w�]�g�  \B��AL1Z�u��(U:?zF����V�I�˖ Z�ʶ�e�Sj��9����A���5 ���x�S���\�8pgTeM묦MKgz��Q@�~ʃ N� �55L��S�Q��� �`� ��GR�n��wIʇ���� (�n�X-�Y�*�*�Y� �bA�%j � V  ȵ �H!��j <�W�"|�0���Q�Q��ۺ" @�z8�K�� �5)3��  �� �~�T�C�CQ
��lƟ柠�� �T��li����)�������� �_- �I8��!c  ���^S-k�����%j l   �ܸ �Y� v3�nUZ+pi � ��V `Ő����u��	DtNI�K��'�`��0~[ ��Y �|���  f}z����c��9s�4�$Ԅӊ�<� ��� ��#�����4h�@�4H�2L��~1 ؿy% ��&� �Q_8 � � : �. ��fDځ �䩓A- �� ��^�� K @�7��q1 �0�8��N��Jw�]���]�z9  �׊� s �N���4�W�1�� � @���� ���G�<�d�ZО�]���U:  ��)7�k r�ĕ ���X�����]- x�� P���
���_F ��5 �3 �Ư���S��ٌ������,�f� (�)͕{���=>��β�eo�L�T����`�h �5�DB��eg�F��|�� g�`�V�J @�(�}
6��7VʪΗ��	��4�ZB<^ }  ����m� f� � 言� t���@��!i^I�_3&���; ��t�	x5S�÷�	 ����X
 ����� X�p�e
dZ `x�����(�ytdƈ����G�*���`��R ��AܹOs���~
�*@����P ���?U �����R�{P3�������M�Q5����҂�+��  �bfԉ��T�~ SQ�iT��m+Rn�6}c��\s�G�
�^W�T�c��)�'�Â��mRK�ԕkW
�AU�hK����!�� ��B/ �A� ���-r��x�������1?S� b���N �8� �D�V�o#X�I�b;?�>]�O'�ى���f�VƟ �c��a��b��~����{�����? �!ùS�( <� �.�ߴ��t���҆QБjx}�
�@�kɂ1���� D��!�o�j  ����}�m\ �A0J�_ ��� �E�i��\��N�2� �0�8����� �H�z� ��cZ��^;*( `�u��+ 0B 4,#ȧ�c�8 0)�\�2���q�~R6f  �_�0	 h��Vю``|g�v�(0�X.��X �n
Y@�?-���SW �@��� �-��빁��	ҙ0y�l.�ih�v�Ss�M-�� f�@ �m��E ���hS�����!?o��;� �7 �  ��q\ :,p�{y���0 ��5�l�*� Fbj6H#�� ��m�T7�{6  �� b� �� �|��y�t!�y.�jf$��M ]�{ ������A  �=�
n6���1VL��|�(�y���΍��W�W���������q����Jli!�4k. (�5�(pC@�2L�6� 8�>��V���B �U�O��}�������(�* �*��K	 Z���`��Z���X� И�U#���C<w�� � �7���[ `)��b����6��� 0 �w:�[�ld�6���\��4 X= :#�k p	� ��^��7���濻E������*ɸ>:�Z2_͔�,;��j-�G�~�W�7�^<K���i��M�MF�G�+w`��%U�_�ʷK�¯��};��
�#p�%��wJg�.y�/�( ��; ���Q 3��  3~������'0����x=����­�� I ![l-��9n�=�=0����?������
 `ٿ  u�7�M<+1�U�R�"�^�/�?���0�8�r���aV�k����4 )�����XG ]=*u+�ˁ�[x|��   дbDZxO��1���.d7���|Lz+�e�z��   �> ��5)]�� �x�.ӪK��ҭ����b��]H��9�IS�l�S[� ��N� ��dBi�)����0��
z���1�[����]Vb.k��-Q1hZm�a�k�k�ڄ��:�\�� [ `�<`�`mel[�� ��@�`��S�c �N�i �m�H�zLN���,w�K�C���th`[�e�v@' $�5L�� ��N�*�:�Q��5�0��j������c�[ʷp��!i�"���J �|�"u���= Ԭ 	Xh���r�����f��:P���E�6Ҹ>�CkȬF*�$���V;ƞ]�S鶌�J��b ��{%  �*�a����@! ��ѫ�����&?���0�� ���� L����OkF�8�f�
�Qզ ��M��m �]F�+n���[�6�l?�_���  ��-7�U. �}�}jt����7�o˹�J! H�"Ω"�9�e�"�KH�_��,�E�p����J6b����k60+s �{ׯ��i�!nD��ؾ K�� 5 d��������= _��<������?-���\v$��~RdD�
� @C�N2
7����Uy����Y`+ Ѐ�7`�u�f��xSo��>If�`�Ä�8斢Y���9�����O}K�7�i'���~�?��1� ��[�9_��� �K  ���~��!�bHq��d�.��,o$W ZаL���eը�����q��waZ�S/����I٠  �c��5:� �5 W ��� ���2< Ċ�x0  ^AvY���T�i�N^Z�t. �u��@��h�]m��	��� @W�TH��I��)4�l��7Kk�~s�� ������s���*�&��"��/��
X
 ���U� 8���U8 h�D�؂ mPP��V!����Ef�M
  %Ĕ��  n�\L?�����z^n �!@�� �	/�y �Z��Z��UN ��~ӱ���?��y��Q�]�/ �� ��z�  ��S`��s��n�v�&�>����_�s��/�գ�#�>�S	�O��]*vā2������>�6�> ��wHOŝ�[q�|p���A�} m� `[��\�U��фt��H'ǡ��ƙ"��&���LG�������������ԯ��JF�ʟ4��R �{I � z �a X���] Vf ���кvL:r&����$ w��謀���v�@�߇���
 �/ ��3�%�L��)E�z0B���s�q�����K]�B������dsZ��x��g ���@���`�m�)�
�` ��G ��P�Z�&�SK�fi ��� ��;ӳ4v9*�Q����vr�s-� �"��� D0Ũ��Ĵ��R `�K�Ֆ��U ���UEhs���*T:*A���-OZ��_u� ���^·�s�i��ޭ�,a�W3
 �n5���@�J����W�u*��>%� h�\'w.�ڹ׶/�x� @e�99  �� 5�PZ� �r2��3r@K~�LgdkX��u2 K�|22'I����Ț
��y�	`i]
 n V��
щV� �����E}���ؙ� j�M�d"�n�壿�/�9*c�]��mg�p��7~J�+n7+�5V�֪�2�K��)��~,O���征O�����{���'L�?��(�K��}L~ lO�_��	�=��g�����g�'��=,}ۥ�`
  H�OI[����S�/���?-�e�Ё���?�N�W}�c�`��g� ��r��͵ `Y�1�7-��

��� �)����Q2G!`� Ffo��	�K @ݭ�R�U���� ���-kƥm݄�
G�V7�}�0��t�? l۫&����4�T��B �1�� -�頠 ��9�� �B�@��@e@,�s �	�I�+^>�ُ�k 8U���6@!@Z;� `��1�j� ��jץ�� X���	蘆�	N �Z�8�'J�� ��������3�- ��� ���{��V� �5 
 �e�b`�Řc�f ��s�D��*�"�����
 �u ��8@k . �"���� @����Z5�����  1EM�V���&�k���9 � `��2�s���oj�� �SXd��l0𕎈_������ �U@@�ݵ�[ l%<d� Z%��Vu �@ ׫�kI ���� ���z����r���ڞ��2� &HK�e��o��S`) ��_Z^/]%d�zH6�Fds�lb;P3,�%��v}��k pz� ���lM�O�����'&�$�U{䣳�̄>�~H�*n#8�F��Kz����w|Y~q��̻^��=�����wn��l��O>9sV~ ���eO�G ���Kv��F>/�8��O~KN�������ȗ����i(������i��ޓ�sw�|T6��)��=!?>�i�@�}^  p�&�2�� d9��� @�	`I ���U�ҺvB�r1� �h\�0�]A�^#��BA���������� ��� ���Z�b����,M 碆�P��\! ���\�N 0��j��0��} �|�s� 23f @;�z ����s�ny-��GL�K� dT��QF�3�44p.��L� *��댐i� 5�Gj�^���ȦK���RM 1 ��	P'�[�	��N�2��tH���p9e�����آ�4 ϺW <��l���ma���6_5 �9F�-:!Q=�:q�L|U�Z��j�� �K�	��;^�K�� ��� ^w5 �ͬ� �����'~/yH6�Ϳo����o{X:��0���t�]�ߏ�Vμ�i��Wv'? _����~-�zX>���N � �����о����/��Fν�y��-[
��ɻ�����.�3}� �n�?��������ކ�I��{�cG��_c��W
 ���@�5
o].s�Z�� �VZ К�c�_���̺�z��Ǥ�ԕ;ɠ;0�+ L( 48��"S����9 ����!̟�R3�΍��o�c�+hs���� 4����� �J�eo�i �  fH��a�� C`�W �� �W�( H7�1  ��"! ��om ��٧M�~l��� Z>��(�r�A@�%�׿�Ē��m�W
 I{Jh��+ ��W3����K�k1 ��3���"Y�,	 �~  ��B h :$�� �$Z�m  T��vp�v�{ ��� 'd���5g� j�iy�  <�G��^Lޫ͌�7]z=��2�P ^�� /�f��j�
� ����U���*�L���`>�<��� �@��MC�e��0k���=��dW����{����;�#_45 �{H�j���;��z������7x��U�K&ß��?���㿑����' �����.���!�'D���������� *�Kw�v*�+�����w��tk�-  �m���99z�� ؑ|@z�w&�/���t��h'Ma�&��|���m�` P��Z ��~ �@�pB� �܍����H ���< �5l��S+�z���2޷H�A��i^M6
4��K��O�怎"�I�3��,���
ޣ�_<��=%��,�l���^؄�l�HN���_��Ӓ	"v@�Pmy�)�¨�1��E��O� �UxZ�)�l�|&��)�<Α L��f�.ΉB�&Z=�k\C��됽 �˱ ��5 i p��#CZ������ŏ	�6�6X4�$ h�r3�,����ا� Z  ��^6�nE��ۊ9�`��@֔4pMt!�G� �E� Ċ /  ����@N/F�#�u�f�cjct�F]�Y�o�u)� ��o�� �U�> �i�c@��-�0�\{1��/��!p�S����@�I� �l�jD�_�/3Jr?�(;ڹU[�����f�Cl�e�ۉ-��9_i��\ 
�|s���$�k��}�,�W��B ]�W�8�z=U> @�C�.-��!�������z�8�����^�^~`ҩ���J���nI��HJW��:w��{�W\��銁	W� ��Tp-�:��S! ��
H:r;�qq5��j �F;b�f� �V�j���U���l�*���N�Sj�٤���K3~'T8e� .���|GA��ߵ�w�9'I��<� �5 �����3"��|^z��w~^�k"����  Z���p�Jo���Ż��<�;9��gds������L�#'�������o����;	�{eO�{D ��}��g��l�t�͕���}E~s�w����K��1 ��� ���#=�;��_�_��5 ��U � hZ;*-9�԰�9� k�1���Q��t D�%:���W
 �Z'�b@qL�J������@�s� h�@ �]��@� 
�;Z�\ �	0 �d�6 8Ϳ��{���=q�!��\H��� @��e��5*@!�̓록Cy���l2��s�b(�7,I�٢�( h�=' �[2�l�9 @0��B����/-�!��Y�m�z�8�] � ��� ��v �� \l�F�� ��$�L��G*��KB%�(�4�4 ����j�j 0a�
 ��Y�]&�_�t�tJ�l��f��� �� �+�JK�� h����4f��M�15 ��wX:������6���7��A2��>'@�S2�Gz+��f������MS�F��N�Q�Nӷ��;KO)�_�]6�}���c���|H:�	�&���쿫`���Q�0z�t�n��m��������]� ���u`׽����{/�AK�+�
��,Y�%��!q�NÌM!i
i��)��6mo�{�z�ĉ���|���=���e�N'n?������y>�̙3�'CNlD/%�7g#�)�PhI�b�C��!�`�J�ܤE��9?w�����Nx/@N��)�fh�E��� C�/�	��MRӫcM�&�r"pMD�
З�R�=k�r�W���@w<��вi��V ��5�5��ڿ�,(# ����)��/TI�:��p�_F�O���՜�Z�B��ע�t�>�@ ���n�p���X��[����������Ju�JTIGR�n+- Bc)E�|)Z�" ��q
�%]UK( �֌���B5�S�m\9���Z��h�s��q{�p��&���0�4�i
@8=*�T��d��r�x��N+�8��� L% O�>>��O�S ��z� L�� � � �Q ��u�;��߄[�>�����0� �Eb(x ��ٯ���a�c����?���#/��B�qC�C��k���T:�܃��=f��������9��v���%��Y@䱐-`�q���wa�h�}�+8���X_M�(�w/��jE8� �����kʑ|E�iJ $�ե�6��,@3)DK@B��F�� ��ɠW���J ߟ��Rz��\J@�����܎C�A� S�/݄>�ÿ�V�,$�HEҔ+� �3��X[VP��UHD-��n��5�o4�M��@��;�	Q|�\��
N�wW��� ���6�I�y��� Ķ Td�)	�~ a��J�6)��P7@:��H�͔#};���A������&� ��W=ؽ)�ҷd�C�j���ߐ?�@�߂5����%m���V ����Z�LEL� - ��3�yL�і � n�\n�<�8e� u�@� (R�.s�J�ɪH@��� �L�q:��x\J˜! ����>���v�3�߭ �]�w~�d��#d_�%e�����m0��7�� �<4��@����S3N�+��,TS���Ah� 4��$  #�yL����J�`ϖ��OƬ�W2�5U�6�ҟ�D�s �D�D��@S?�X�+ >y�@NƁ�����7/�&�7�汧�?P �X- C�~������wKB��<| /�������ױ��L�nb-�0FK���8��?H`�!��|�}�Oq�u�3�Ѣ������ܡ:��P��;1�݉o�g	���Q��Ɲc��;?>A�����Z T�t����]��&�����R��=��(� Q�>�K���vC ����1��l���) q40x���( �*�� )�kV����%������`�P�p�� r
@u���9p���3j3�:c���	�V �%��S���H�*5�����@K�� �A[���`	��L����OW d�? �[h$�D����ZnW��萯��%�5~5x�t��1!�����؇��`��e�P��\&0�V? ����E$��j�脼��Y��Z�Lu"l	,E�_>o	�ǣ�B��v2�R�g�ZĆ�ə�Y�7�v�΅N|$ 	��
�!
������_ǲ�[pt�	���37Á#J �8oo`9�^��aS����]�`���r��X��e0�H	k������a|��7�Ϋ�o�w0ΐ�+܉���љ���ɂ�5���H	��Wq��Bʿ��>��o��X�S �3��%�_� t���,�.�C	��g�p����gA�� z��<+��g ���lc���`�w��g�_:�T�`<[ �o"7�i.�>��t@���Q�c]`��?�P�fA�V"�[b[DXۗ�9���Uj�A�������Z��) і �r*	����)������ H_��>A���:d�'�<��яf�*�#ݏ��&�1�m	��r=�Z��G[��H�h	��O�RtU-� ,W#�H��A��~J@�|�F� �����nc��a�kу@zw�w+ ��o���]��.���3���a-�M	��N$�~"]��I�Wx�r����� d-Z$���� 7�H���)���~�}�C�_���YL���[����AJ@`/z{��g���|��l/�W܊���K�x�$�v돱��&,f�K���*�a�����t��m,���@�vt���F�󷢳����������w~�r��CE�q��S��XR�G�(��K���r�.ϱ��H!�iga��i�4�Ӣ+��O��3�� �~ d������V� 0��6Q 8e�w��w��
G�\"(��`-^�K�T�k�:���Qw	`�)�%UrnV�U�������,�[��R�s�k���C*��,$�BC��P�V����P-����R����fe�zK�M}% ��[~���g{�`h5L�H%C��렊����!�m'} d$���h��q��Q d��R��K�Uӊ�1��8��A._��$ �I9Ù ���R ����rV�����Z���r�~J����0��������%���.����.]��71`D�����G긜U\�KP�a��al��o��oBK>���^$�� B �9��E j(gU,8+)l�׸<V(!��O�W}�g	a��Gh����u�L	h�[�cq5�)��v�QxLus����O$�Ӂ�-	`���������P1�a�6��V
�7ÿ��o'i�1,�U�CF���
~R�uk]���<���ÅSa�*Xa�m��!�����E*���*n���q3��+���IN�)�r �mT1n_����n
@W���� �S Z\�>�a��(��KP]�r�ǎ��s�Y��� �B"6a% �TJ��&F�]"v���睅!�e�����\Q�q_��s?՜��ιh!P �( I��J �, N$�p�- �" �|J ����΃N@�P�h#�;���=��w�[ ��U��=2�5,���w��o�&�) r��~;�{�{�O}{Y`���ڪ[��M�᝟�7�~K��a��VU���C��ۯ�����"�c����!����5܎|��,lY�_\��{�5�Ipi��p�u	�'' Wtp^% �Y�%�z��f� P2�΁iW�tE|r �m�c� �o7=��@K����6򸛯wQ �3�� ��~��9PZ zDl�������Fl��@���%0�

�}��� �9G�y	��&e�K $���3
@!בwT5s��) ,�:B�������۫�����Jn���`��Z
\��R	�t��r��@�sZ�M��{��������r�~�:��6�
 �K� �-A.�.�>� 'h'2�Us�;Q���1hj�|B��b�*�-	P�+-c�uOp�	�� ��<��?� ?C���T��f���|�:i"���~�M�9w`%�(�2���ѕ/�[V� " ��a�f1@F�dy$-"=��H�TTx����"�����H���q	�Sd٨	��-E���z*��0�`���@�- �y�5HIs��Q�(��?� ,��R�J � ����b ��ܯ�P L̖�)�Ǹ� �8����/ Q��M�͏�!�q*�K@n��[	'�q ��Ϻm�c����a�'~<w����A�aJ eA	�>u:�߷C~4`���G(���7N�{���ϟ�=N�<���@(����V,�EXH'k�R(���͗�o�}�r����m�c���p���w' �s& ��Plzr�gk�"�	P"����J�M�a!�ǚו�,�.-�e�����z�Y�f7�(�Z�(����o���/ r�Ycÿ�5ZLu��
tT�f�S��YK�!5���fx��� 4P j�ע:��{Y� sJ	���f֪��v������uūXs[M�LC $ĥ9ߒ i	8=h�2��RZ���ҡNj��59KQ-��cn+�k����9��䎩���Kd*�s:��ڿ�~YZhd;9	�u	���|�k�.
�-�JUS����Jh'����<n?�O�o�># �
��E��e;�j�1- S@3�Cn�nM�TP5ש��(aO��g����Sn4>���q�)=��%q�Wp�VȔ2P�u]-� �qԗPʸ^�?��mB�&!�q[X8�Y�T�'ÿ#d!���?w�O��O8a�E(M�]�s&`='�NLG ��G��N,��;� ����p�{�+��N:JX� t�^��2��t�z����6���P/��n�F�@������} �X8��s?������׏�׎�/?|�l�F1�v1���P�&�m	f9����w`�`/F�����~��~pKK���w-���8��~�	�\��X�9�j�^
@��-� -" ��/���V�L./��ЕC	���}{�٤��w� ��]�v�j���s��QG��o��` LC th�� H�t�jJs�JtT�f�S j���O։pJh���]_�A	@Ukx" ��/��PA���� �1k��
i�-X�Fq�)^�B{�J"eqP�}��
�x�"�^ �D��EŤ6w��a"�"�/
J���S"��z��0��%@K�LU��9- �b�k�g, r�+G��SV��H+i�t2d������ �
�@N$�
`���o#��{I��TИ�&V �ݕq��	r��`�.�0�����>EP�� 
@�wu��/[�F�?�i���Bh� �U�%~���d�߮�K�KKX[��o9eb��L����%�,�>�O���~ �"��0]0/�H ��i��D��'38% �@^� 䱐�%@d�� M�N�N���]zz�v��C���8N�ܵ�{X�?���O�
��}����*;�R���_��mFJo�0nlw�<��u�aI�A,.د��E $��%���;W����N5��������s˽" �p�������h��,@$�E&c��t2Ҵ� k㴹pm� ��j2�cf,� ����v&r?�� �(�d��t:`cK����.��a��Z��mP� ��
`��mߙ��5hw�DK�2.3k1YK(3�t�:�cpS 4��cO4�����s[ dXZu��Z[9k��6i��\��j.O-���Fh��~)"PC�܊��41��c���"�����0�A�%`� T�O�Z��.Z��?V/�d?oڵh.��(`�˝ 9o�N�F4��j�6� ���{����B�z���/�J��{c[ ���e�/����Q��D��+�Ϩ�.��Z�DB\:g����?�t@<:�u�_�|�v3����j�k[���\V�/Ҝ��$�@�ۉZ dEZ�[ �
7��+9�;��+����n
�U��W`~<��=�T�� ��NU ����US4�ڹnX�Z�_�����A���?���V���
���@c�2�K�WZX�P��u@�� Kbߧ	�F%`r�OF�΃�E��	�`"�o"�|A&�B�% ͬy��A�d�H{�H�P��;�wP v���z% ����!|�Y�,����'��O�/����oVw�[\~C>�y���Y�ť2��a��J�p�!�\���P�*܍���(�AX�`�KG���]�#r��P�n��x�>���O��o��e��0�B��5_���;�т],��ڿ� ��y�@:J �B����߮$�kzrXP�נõ����h�G��6����@P�Y X��	ƅƩ�
��|�¬�����\��¯Zj�" �N�����v�nC[ ����f
�u
�Y XK���,�ظ�u K ���R
 V�r
�

��3 ���H�@ClZ�!�@z��s�����/��+]" �
���>Ta��t����2Vz�H��2E	�S���F���^��涋G�#$�	
�2
�

���} � ��L�H? �> S	��}�*�g�ԥ�U�¨�r��`�z9�	��^+�@���\�A�:� 9P<�:�tC���)� ��`>�}J�"���>�/��j�s�rK (����& �a�χB �$���Q8_����:�}�"�l�B�9�\T- ��6
@;��H��
�)è�- <(;ypv{w�p�Q5������<���XVv{۞ı7����*67ݏ�����������j���ڻ������U
kk�Ī�;���l���*cu�(VW܊U�[�&|քau� ���X��ӛ�6tևnņН�R}'�x�7��׏ai���V<��x���0���1�5�+ !�i���@�0�{;�N��.��=2l*�G��YH2L��{) }`Ȼl��
;��@^�+ z�������%PD�/��r�zE�G���͚w��eh�`!F��KFU�g��W",p*�x�� 4�W�x�+ �>$�IcKB*�r��p��(F!~��Z.S=�E	�F�s���g�_�V����ѿ����r=V��`L������6��Z5kqU���@h����%�e�"�}����%���_��v+� W�Q ���H�#]s]����S�e�aШ�?�7�0���Z_m!7I�V ׵H�)*��t�~�=d��{U�k���� d�<�DH?
�0A`hEZ � X�Z`]pf��:.(�A� �G�����F���\+QM*)"a.K0W��y.��mQ��eI�rJ�dF��:��� ����T@���BiX�}�j�+崌�嶁���Z�	�Y�W5��o��/�>Z"�*�~�T� ��
�I���a�@���_�@��*3�$�&�-�#��Џ z����@�� H��!��T�C�'R#,�XZɔ��O0���O��5~�~�']��A:�y�v��� �f`{;*M�����.������x�cw�=x�'�Ě�`Y�!lmy���cx��c��o�/��L����.�>�������G����Q�����#ߍC>S>[�y�|���O8��w�_�3�^�^$Om��z�,f!�Ț�>���&� �^�����#} B�����uv+@3�V��:Yu����]͐_�j��,Ԭ^�$wKr-����������TA�ʲ;�����j �6�r%@�̤�M	p�Cg�td�Dk�r4�/� ,A=_m�b:Nu�c��d�g��{�!�ͱ je�_c }�C�Ij�y���:�)Fr�Ԫ����a�s�X�7r�� t�3D) ]u[) [�R�	�,`�A_��ҳ���3׹u�(B%L��W�P j��QW��E���eA[���/��SKZ˹�K��)-���{޷}�;}�[� 	�>�*�H�@��}�_@� ��-e<	g�rq�d9���,��&�� 5{����_�k����Ct�E��b2���xT�?CZT���p4�f��,KD T+�jXC^G[� LF�`{S�Y������@Z+�ղ���ƜUh`�ב��=��KYS�`X�+�<�|���~ר�0��N��L� �G�����uK����}K��K���l��:��IC^]!`#�D�׬;
j���D�\a �D2�=�}��" \׀ ?e\(�聏��6N"�`��D[(q�9a�d���O��#�
�j�*�뚚�(�����z��7��Oem?��zA�.t�.�E���$Y�#��:h�]��m�F(t��N�5� � ��_�Z��������2��T��xw�~wO|�-{��
^�"^G6~�l��L�|�m���"���5|�F�~z�W�Ԗ������_�{��/��_��k���W?��W}��xw/�n_���O�P�b��d'>��%�����0��|�'Z�N��9�f۔+�) y� �� MY�ha�����˳������^���Z}u�~���T����  ���Ϫ TISk	"���4|�ev�Y�N
@'���Z ��1��#�H�tl�:��P�Z�H@�*4�K_ �@���q��p�3��V�rݾ�^�� ���z�{� -f�?3�������9 ��V Ʀ- ���X z<�D���j�e�[ $�[Xn5�F���г��0�2T���gm?�b�g�1�	�_&k�<&5�����>�~.!,a\��}˖ i��*ᶴ%@S'-{MC��.��sR��_DBa��|�|����a s(b�n�r��� H��H��I�_�Ͱw#��qa�g�*�/.B�U ��,ls �{[�.����S����A)t� -��n�}�M|��7���&Ja��,�݁�����D��#���܊1�-��V,��Ln"G�B�Q��H�A��W˴К
�D)����/��ӭ-݅�?���g�9��Iг����*v��a�©t�J���� s-��v�B:X;��z����|u�ٽ�I"��ah@��	���P��L`���� (( � 	�*W���J��\/��'��m�:�u5@��fXy��[KW��l%����h.�/!�����������ދ �&�ED ���N�/�M�ڣ�Y Ϯ ���}� ���Ȁ�� Q����+ ����𗲨�ǋ���E���
@�{�U��� ��"�=�`�ß�D$�3FP�}��ǫ�㺍���:��>m����,V��º@K@M�*�YS�^�%�i�\! H��x���B����h��7k�01oS,��K�}�Bu��) f��ȀY��?�B��.d^���/`�3�/*��b/<�x�{i)J��A/������$���b�+����Y��p핛����h�n|n��Ե�/~:ƞ�qc����>쬹;���OaK�X_s;�Uߦ ZCVW܌U7Y���Grc ���A��Ǌ �te� V�r�C|�~�Q~�Ql���o���;���6��/���y�>����fص1�cj����D�|E\��ru�l����R�t� �P��B3���D	h�^�v�RJ�
tzVS�֢�&��+� ���X��$@�m#��)� 8��� 	�����\��-s��И1f��S{�% U,P��z
���@c�@� �� �vֆ:���
tU14�)F�X5�����f����F[ ֳp\����`�O]7/���@�@U��:N T+@Ɋh*Y�&/a�7�{(�D����!���5@c�D 
�o��?Ë`��?Y $��Le- f�k
 �.�2� ����`w8l��q�lJ��]((���7[7�@	`�_�/5V6���rH*&rzRj�Z ��u% - ��13�0 Gc�g,&�� ��_����S����DD t�����B�E���`"=�k�3�i"��|���Z D:�S _f/C{`���S�O� ���� �I�Έ~3���F�c��2���� ��Z��I�{��p��ﹸ9�� �2�/���r?ʮ�GM�?o���^�6�1��X�$�4r�]� �1�Ե�����²�}��~������x����描�/�o�ϯ��?��&�����O�F�����
��O��/��#��?��'����������E��#~�+o�/���7_9��_9��p_��m*;XxlfME
��/��h��7y���Pj��©��V���g��ד�0��z� ���# j, ���BR5�[�;�:�P�*���F���&" V�k	�)rc��Fu5�}��1���U/��
���5�t�# ��lD�n�ⶫ؈��߿��%k�W�����4���U�ǂ���-S��Y;��X�6z�EkT�70�d�7���5���֒ S4f�_��=���i���� X YП����@�5"� % J C_#W�H�95�*!<n;��¬��y�4�W*�u-W���Y���� � ��7	��>	fG�gJ+ �}DNp_�- �TQl+�_W0�+�&U2��)	jjS����OSU �ca��u�ǟ���R�������>�y�eǜ��� N! )�L�S��������E��{������0J��d�W!0��y����]��B뜛y 
�+�;�Ē�[�AI@�6,�ހۇ×o|߿�g���īw����K�~�/��~���5^y��x����^�7��c�I�m��Q���6x��?����z��������w�?����?�wn�)^��U|��o�H��\��,�7��ڄf f�7��A�9��FN���p�`���ZI	X�z�w{�+	�}	iM��Н��.��9 �u�=���?�Z6�,|���H$ "	`��4�9-�?��bJ@�$W�@Gx:)���^��U,��wK��z��ס�|-j�2����� �0ehI+�� %Ŭ��P��� ����*���N)r�n���OP(�"ZD4f�_��t2%My�r��������xX�s8�Wu|�$ �HgX	c�?���NYn��1)�;�.
����e��/��g�l
������@9Fc>/hp� ���� ;�Z{�p��<�k!J�5�3�w�Fz�k�Z� �
��/ њ��o� T�<�T�|	s���,a8�`6`>`��IH�8k��d�K��T�~<��c���s��Od"��Ⱥ���Oz�0�
๤9�� ��2^��j����T]ۆ�YCXR���;������{�m�lS��63���ܨ�����t\���>���l�)|��m)����1Z�����~����XVӝ�
vl'�LQmT+�dd\�����dm�M������M�~�E�1��Gj~�,Ԓ�(���<(Ik�,HT })����!Գ�i " �,�ڲ��=�A�bйX�u�SЭ֩�^�ܿ{��W^.����l��8�����S 49["�r[���~�7W,(k=�2`��`�}
`��2��a��.����6��/����(D,�$�m̖S��!�bֈG�"� �I��� �?����Zɐ�Zÿ���k�L��kX�_���U���j����~6Tu�|�US0ϝK�US<�@�ɷ�V9�Z_��5~�E�����2 ��չz><r��!.��;�O���ԝ�H��%��&%���F���o`��3����u�F[��Sk�p��ׁ�1@��Q�B��&� �T�Dߩ�_˅��% ��OG�H�\	������5�]g�r
�J
�%݅ܿ)Br-�4�+�y��9~���GZ����cA�)�`U�9<�E�Y�o��/��eh�	CV�(��f���q�q:	���~� �+�n��%�J��ǀ��	s�� ��� >�`��&L*�>���_�$ �{���L����.�K�	�)0E!��a~�F.8��d�π��X�(j�wQ�D�E��u~	�왘?c>P R�i� �|<��Ǡ�?�YȖ��.��}A.< ��b�2��X[-�2��k��g�W�iC��n��_��+1����7aU��)�	�J�b�{#��z��N%Cv���"�{�[B`���ǃV�˰��q@���f�����c�`�n����l��8�HkNHg?�������&N�o��( u,ܒ��b�en
@����S5(�4@
:KXH�%ԭ��'* V��d�6�0�P�$����#�, �lXb C}� hN- &�j ��Kk ��\(�<�.��/CK�!Z��g�;�
�An� ~�*ԕ�@u�rT���,�e���IB����20�Fu��`B��&��D����X�,� ,G�H�����C�)ɭp5��L��'-���h��s}pYX�7�T�y	@�g�H�	P�s�
@k�rK�Q�[_ˠW]j�+
R�"r�}W�훨Ӌ6*�71����c���&������e�W��N :� H�O��3މ��u� F�*�m$����[�/�O���o�� ��G"� �a?�Z �X0I �) V��"���3�3>)���w+�\���/B����_^��+��J�c�v;�3u��k�ڻK��bK���x wb���)?��0�חxY[/ޅ�E;0H����/}䴀�nZ�@7k��'�~�Nt2��~C\�]#��֑67ZX`��7����9��k@+���N� tR ���[��ﲂ~�`�H�s2�{% 1�թ��Z�XP61TJ�K�D�|�(�X�M>o�rԗ,Gm1k},�:�t^)C�f�A
� �))�)"� ����3�Y+��n�+����}���K��^��i9�19���G	��g#���4�>$����^|_��,	�1��763�u��!n���@�O�n��� �fY� �5 V ������g�zٙ/��Vk��3Š�
���r���/�	�z���)��N�@��%�b:��p�OHǈ �g	����/������M"H�|_��	 �]�ޱ� ��W����p�B,�h�
�� �T��g���L�_����#����.�G�%E(����ޫC�_W��Y�he��7e9F7�?�߿�/8���܅=��qC�#�U� v�����XUvKK�a��F��܀!�.�T�nG_k����G��h�����vui��<��B�9ǧi��D�p���m�ʿ�Pp">�5��%�9�5|����+,(Mo�A �U���,*)�1������q���jeA��� #�7��b[ � $�
qM�hL��/���_�E�2�1c4� ��:��A.$ 3�MT�����)� �h,^�F�jP�L�.U��5x'P[8���1���0����*�5,���ׅ�l:(%8�(�yc�N8"�2J_-�ZB��EY �"�&�_���Ǡ"͹+Vr9u��w���|V�k	��{���}���v���$�Xg��%�M����Y.�#�d�� S :�s��S%�P�)�vB�u
ϖ������X���������3�A�9hA>�p1ԝ�	}�39�/ a���!� �ޗ3�< z~A�`�� X�PK�S�Z
a/ć��<�`"�����_��צ k_�};* f+�Q}^v���.�~��( �\��/�E����{QtE9�WPvm%*f��qn/z-�X�&��كO�{�O��~�x`�8z
��ц�c�S�~[�wam�f��ܷ�t�~������z��/7�&�� 0��s�������ÐӨܦ���i�;�EXC3�4�:�(M�	x�p�@�={�c'@S T�?U�7k���
@"�@���ߙ��W�\���� ��3 3��X@i�����(z~%,�ԕ,0Xkj(�Z������=�Zu�cͿ��Y%��1�g<VC�9[�Z�����;�IG�~�v�M=�e�HBݪ�s������e�L����Ϥ �R j]R��
�����0�o�~��
���C�� :E �<#d	#h&r��v��r��vCV�(�1��O	д殍 �߬�]z�[�z�g�
� csX�s��i�3	�=W�B���Q��ڿ��rπ"" �W����&�=�~	a��7qr'|���^�����" 	Z � ��n����sU���_�C�5��ϨA͜v����8u-Vyn����K���u'�>���џ�ٱ����/�Φp{ӗp���P�06W~
k��a,ĸ-#^�@�ܤG��N����H Ç�.ȥn9�ך�%Gpa�:�5��'
C]�\mY�j�Pu�>O8	~�_S �2@�
@]8� Hs=��+ �V?t�w����X����3&�X �`7��q�EUV�G@#,L���,D�XHZ7�Z��֥�;k����=)4�0
d��j� ��װV�}�~��)�&�B��@�� ��X���3����_�S���$gK ��)$
��
�I���PG��"��Q��H�ȸ�v��S\���V�m9+���M4MR���:�o]�'�o
@$�Ӭ��� �� e6��7`��>�"� �,p^�)��7P�c�|�_����LG ���S:"8�/|$ g�XH�x&�?�E�s�������eJ�����ld���RM�yȽ���0�/+G�A�_S������BW�8�3�bs�M8R�8^��*N;��'������x_��
j�>l�&���5>��uOcK�=XWyV�o�2�����%{(�1X�E;�_�}�[Uo^�nWֱ݆`k�|�~���'����-EM3kȚ&w#C3�H�E��	��Չ��%�$^ � ��> �{1�7��U R��܉Y�TP��g!$�� ���o��t�7u�P��P(ab���N���ÐwoB�:�/�@6�g#��NH�^ӕ!����8m�`�L�\�V���3%�Y��𧼨���<XkH-���Lbx4�M�`� Te�D�VH� ���u�!C������@�w�tR 
���u��N� 1�����9�e�Ղ�k����(�|,��������U�g�-��|��gA�敩`IE��Y>��o%R:�� ����
	��q��X(z���}j�5�|�������QO��\G��f�8�LR�[x<Z,�s����[y,
m<��t���дH��t���H��s��_���_�%���6#� �?�KK�-Ε ��� ����D��V�[� �����z,�����R������5�=~G�߫�RȐڿ��7�s���Q$x-�0��Pb��(Q�"8��/ &�8�Ba.�Ae��0�~���ƺ�}���p?�V����+ *��>�S��o	@&��^�V���_.��\T�z�\R����]U��5���Պ����I]�e�7`g�]���,���g��'p'q��7�_��om�=��6l�:�mG���u�ck�}�X-��`E���b�lFK�`�t7�ף��P������t�O�=�;=ր�<����DVEha�k&@�$N8���, B"P���3\@�@*J�F�r�Z"5�XXBG�.֊�sV� ��$-yʶj퓑�_�+��
|M�J��W(�3Y�ڴf�p�Z���14d�@���R�Ǜiuz��
�^��&� 1��_6r�/MLHM�|�w�u'$�u�b��]�s��X������ ��{2ә')����|O� X�"�S�V�k�& ]Cӈ��5� �+�ܚ8�(��h+]�AC6ŝ4�ؕ�ZN��zDN�ht�
A.���0j�������DxO���\1p��5����Lv+A�yb��I��W#���[@l�[ a{*��(� � �_���T0鮁\�

@%����c�<v���Ǡu�,�H ��#��"�]�Ek�eW��U_׈�9hI� k}�s�aO����|��_2��
��?�9��������7x���x��Gx�����%�m�v�=�͕wc]�v�ނ��#�(?���}X\z#�Jn��w��[�ﶮ�Ot�f�A���c��.����7� T*	`��d�S z4@�3`�{��}9dX�~wk@�C ׇ\�(H	��Kj��j�Yu��L~��}�s��V0�F��\N ���ܖ�2����[�F��'��1��s/ �9ހ�����&�z�s% �<����Ԉ�Ⱥ�0�y�ݤ�A`ux��{Rh̰61@�-(v
��V7�j����r9#��K����G��s�4�V<� �I�w'� X�&�-��s" $�}P#7��m�e�o(�<��G�H F?��V�{�u�_��>�_F��jT�hB��n�-����X�w}���گ��c�	%'��'�)��;x��'�=���<��:��6%�8�(�ö���}�W(>J�� ����H���Ŕ�"J@�U�� ��-� a�E٧ K�SKK �A�`�������3�߾��ed9a({�5�'����XRÏ�3��d3�m$ԝ��}4�ѯ�a/H���q�M#��u\�^�,�p�j"��V0�͠OD|�'�- ��4񅏉�&� ��ic`�Z,V��>\g1�����g�k�J
�_����$ ~~e6����	�X��~�
 ͹�
@��� ��+@#7�2��(%�ϫpw�#������� :�%�#��� �K��W�U���TͰz�w.Z�%Y��9�(����C�����p�O��q�
�&E��o���_��������5��%�븳�k8R�,��<��`c�SX�+�7a���U� � ���r����Q�(�`� l���CK� %� �4O! fA����v�3��Ր��\Z��fE ���=���?��Oo�amg��5��OKθ���;��p[0�FAҴ1�OE{�2uBi�zj��f���	���*�� ��R؛�$B���N�d+���790Cߔ���) 5F�k�@_s"� 2�/�4� �L~��zL�T��ZvD �l�aoc�[�aA�Y��`�]�`!.�Y;���c5D:CꎓJ��d�k԰�6S� ȹ�aE������S%��1�_:���:3C_ցLE����'�+��x>F ܚ ׇ�|�/�m� �9g�0�/� ^�' &���) Z�C?�;��/NH�;Q�� #��1�%Z������������ �+ ���wi1
//C�����u���ц�y�N���k+�ނ���#���R �l��g�3�U;�;���ɷ��$���$�{��١���}?��=?�]-/�h�s���	J���XqV�oÊ�MX��ʸ"r��.%C"�Uru�a[�� �z��\	0����I�o��S
 Cz�%" �(In�?9V �H�K�@- �
 W���y��K�(͔���Y�9�&ួj2|���@��Pw�%K:�M(ZY�֒��$�,�l�],���YK!^� ���ӗ��Y LbC?J|���8���&���&Q�K!�H���R� �}�� ���>3���(Rx���
���B
q�?���CƘ� A]i_A!�����XwK��Z �� "���`�����p6�$:����&�}Cc>O���d�{�;�}	��G�A%����Ϙ� �(ȿ̋�˭������Q�����?�g�{�ގ[C�����՛~���/p\R���� �H��HK�ۿ>�W����>��3<��}���Ui|��Ƕ�{���N�݆�"�1Q�_I�h�n{�W" �
�� i���7F$ ��V���&��C �N��j���x���w+ 2|����]�`��.j�/����d����5���U��QO�od������ZgT ��5rr�$���m��0䄜�ob��`���Gh$�{A�k�R�ZN�w�թ��<C���S��c�E���~M4�u�E�[��D��5���@]��K=��=�H}\�D���71י1r�r5*X��k�D���+fș�o��/�7��ޓ��S	"�},��S��#���rF�̈J�u9����\�0Ex�
@<�p�y�PW����I |�7��9�+g�;-|��?���! ��e�� �&( I/D�'Ґ��L���|"Yj�_k�υ�ȹ����QxY	J.��we�Wף�f��B�j�p����O��g����g��x��~	~���"�j/�#y�M����������g^ã�?�]��Ƒ��cw�}�^{�/`]�V�	܌U�#X^zP��z�K�v��h������r#J@w�5hG�zk ���
�Z�Ր;�	2��9�ZS�r	�hh�a^��OD�:�8��ܵ�4QJ�r֡��=�0�4xS�P��M A8�pj*R{Q�����P���q%���L�Nc���%�m�Y�I}|����t�����<p���0Ĥ榐 ���a=�(��a����_�D<�w��frox- ~ʬ�i�W�rYX2P���@h�H+�d��$-2���u.���`��D���ؠ����9��`���1B� ��3�_�'����AYScحC2�, ��(�}��o�Hhծq���P�}_^��l	P�O!��1��r/E�������%��GН�u�S�u��u9���tB7��Z7��$�D�$�܍P���
�~.��x���y������x!�ha�%|����Œ�xteI��X��ZcfX�f� Zu��[�p�L% R�ϑs�r���Ŭ����
?�WU"tM�:��0��c mVz�`W�ݸ����l��G�� 	}I��,�O	�+J�(������G~����O�� w��@	��4>��5`s�n�ގ��[���(���쇌��K	��\%P�]�\HD@��E������i17SQB�*�%BlMݔ��?N�/� 4�U�\
�u��P�%Jxp	�<дԱ�Q�"5M�tj�LD��f��7fI�=J3k?ND��{2�y4��k2fКal~<�/ ��ob~��,&g" ��;��z�3�tA%���[@|P[��N�/8�j&��p6@����}z�+}�� HK �C����`I�RU��`�ÿ���n@Z T���#�H �LG tӿ���P|Eʮ�u%��6�zf+gw�c�0���=���^�U�,>��
~qӿM) r}�;x[I��|��;8��������C��/��O�����_�і簯�)�z[(�wb��V�(?bK�>%�%�1佞��(}�r��-�t�R
6PD�������D�㭫1�e�0S��p
�)�K ֩��
�~��*����H��gA5�G����!��4���4�@pG�:p���^�1��c���|�>����)�5�/ć����V�$��C�
@�N�/�a5}b�_s6@��%��6˱0�m	��4�g0T�Vd�l��QT��,�H����@��]An��:�q�1;Z�:v]����s��B9	�W>�3'> �iI=Жl�e��- r���r��/ٜʥz��|b� ��m@ͬ64��Fg�(�2�bu�^K ��ó�� W H� ��D�\ 
��o��;�9���;�������o�d��qO�K���y�y;+�܋�"�۰�3��V-2z��B@u���֥���m�*�J�L���	�ҚG	�kИ`������z����Ci�Q0��u�'RP�Ҩ������xD ����vthJ�X�2��?��c�`jd~�f��c��&1�O��T���M��e19WPOs,	�s�&:����ׇ����L���p�H�P}�$�}B�����0B�,���% 󼿉@|�;��I� ��2/٫�*��U���h+����&�c��/w��ē�2@6\?��E3���B�H �������04	���}ʉ ��5S	�I�<��f�;��`�KgS ���<Y ��-���-��҇^ T������� 4��Aע%j�5�����>�=M�����2߉�������ߞ�)_\�<7�%�5���M���e쭥T?�͕�bC�SX���s�!L���B�F%��ף�h��w��B�M!�,	�B	��,�:��κ �W�� h�6*] �]jw*H���P!>���v���i^3h��C0CZ-;��j`�6p�n�\Fa:Kb	��_'��b�Q�o9�@�
Sar�O���ĜEȐK��N{r@�X�,�`�k����ɧ �SN��m"�.���`rӿF�ޡ��8w�oL  ��N��<�fY�s_zo��|
`Px��+�Q~UP� ( ��nG�^t'�a8k���Ǎe�㞚/�َ�
��򜍜 2��DP���8~r�_����g�'(�u~K�	�[�i�y[*��
��Pp�e�1V�W���"0���^[���E$���`��V��_E N�@5��њYxjT!ʃ@(�hpB��3���y-�`u
_!f�X����m�eL�t ����X d�I( �����o�q��� �,`q�Sq��J L	��ҳ_�"���79]0�s���� �a͹ 9��9O@�?�5��O�Gp֙���IH�8	Y�H���YȖK�l\�t�}�� (��^u��
 ����]3�-�ѳhK27`C�>�-����1~yӿ3�U7�80�i	����<2N ��ߜ���/��#>;�<:�=<��2�{��������n�ݩ$`��u:`�� ���>{)�9�z�{w��x�:�c��T����pa���V� �z�䯋ЬN	X4Q4����q"�Fh`�k=�*�Y�-���p�ǓQ�܀����N��4U�e����>P&	 h'�Ќ"��9�E:�i�\�I�ϲ�+��4��85ՙ�\n,���5&r-{��y�з�+Ą�H ��g�&zJ�FX�����Z��}yL"���$ v]J?ݗA��7��LO��@jZN��5���9���22��U�� Dq
x'�pf�P��ඨ������rs{bC���ga
��h$x\�̑�v���L-�	�d�<�
u
�Y �Z �F�;a
@�����o�c��r	�wF�DD�>�c�>�^���+������>�����D	�ukp��A�1��!����F�i^wƔ�(� Ǐ%"�KP�m^��/���qK�+�KXDH� dS �" ��>��'=�\��\u������`� h	@���nNZ�/F_�2�S 6�����po�W�\�� � �O�HC �%?9�����/�|߯�T�k���k���Y�oz
;kĶ*:X.��}7c�t,?`I@��C�z��Āw�}� %@:�1@Z�6-J,�U��&�`vlb�71�OE��F��J	��8��O��i S L	P"`H<��8tH�S�����1����4�bAb!�`�����|�)�ķf$ַ�C	����Z,���#��u��� �����+ `�N�ob���PP�FM+a�O��n=��ؖ 3�c��� �/ ���:@_&脞G�� �� �]d9�?S �^� Sp��O���AD��p����8���N�����c�ds�1�?WL) C 3�-X�� ���A]���`})���ؔ�( �վ�@NXi "ǀ��p?���z���s���#���#���m��c_ݓ���lߋ����.p;V�)��	PW�xw��#`w	h/��� ��l�� &f�L	z'dP"����Ǽ�����Q(4�£����D�<��M�B�*`cv4e��=��:~5�Q�7�>� 8�0� h	����u�\� ��CT}v\4�LO�KG����8�,bj������aO��;1� X�Q�NM���o���ϖﵑQ-	�'����~��|��!���;�T$ �7e���'��M�?�=��K)p},�S{�P$C _���
[ �( =J RW`i�&K �� |�w����?�U@�A�x���$~|�������������^�|��>�ݕ�b;%`S�N%+�7�� �8V�#�7bq�� �Ɯ�� �~ f_ S L���BߔK��& �X�Y��j
��([��H�h��</��,�F�gc���|?CDc����|���@0�)읈#㳜$@��*�p�:	Ɖ�! z ���;��"TN�N#�N�B3]�ǔ ��E@���>�/A8���W��}�
����д�"��U� ���j'�5��L�?[c���eK��������'����� K�p���g,Wܗ��y*L��i�x��+���LG۹�bXC��7�ң��m�ϯ> �P R ���[��@.T������_'�8�����4�{|f�xj�x��۸��P�vW=�m�{�1x�uu %@_ ����⢝�M�Ho�6�l�l!2V��2p�{& n[ �K1����/R- ��N- � `�#FP��C����^ $|e@�~��p�|�kfh�A��N�� h""���:
Z"��h�?^ N'���� 8��/ �S�$�H��B ՜��q��Pz����jp@�0k�&1��!	'�7:-��z19��X�e������wXH��(bO�� ��_��8��T������O% ��:`�
���M	��`s��=�N|��g�/ ��-y�\ mj��ߝ��7�^X�G<��x��U<��M���<5<��Ķ�{�1,}�q(j� ������P�% 2P�@whˍ}3У����B�g�#�*�p�P} ��O�એ%�pQ=J���_0�D:&�r@�%�1�1"���0k��u"� �)-&� �>�3ا���8#+Ձ�-��y	z��
�J�#�|:8��\�T���S��V LɐN�rU�3�@3?���j�7G�S���F�1�52ƿr�@V<1�j`���m.�T���� �B rO �cY��&f9E��ύ��X�{���8??�)���� dK��
}�B+c��� ̶ ���A�����r
@�PE�Q ��0��F( +) �������_�����zE�9�o#o}�Z��`Ao�ߟ�O��^�'<7�s<9�}���5|��K8P'���
k��Ձ[���&�ʀ����-�A�R�@A[(�fu!u!ґk	�\
�ifm=
k�6Mv�7y8UP
l�XS�^�k9w��1
�W�]�΅ �t3�	��oM(U$����w�i^'��$
y+�ϕ ��4��6N�ibI@*3-�T� kgU, �D@���2]��a�Ka��P�:��B�6��]��2���W�F0���
�a�q�dp�H ۡ�H �\rS��y,�`#V�0�;�����3��Z�6J Xx3�^�|]�0�hI�V.U3�K �������Fn�q
A�����4��@�\�&����c}j"�ߣ�����p>??O0%G!��&F Dp�����k�%��h8�u��~i�pbR�ۄ�d8�Ӄ�:!N�[��bM�����<&)Drl��2�O�V��� �O�M�h+�'�M�EX�ԋS������G����w1�s�saÿк��R_�C�U!���E��&���D�~t.X����X�چ��Gp���{_����L[ ��i!P{�`�B??�'|y�W���k�t��p�7qK�s�_�v�<���{�IF��fI@�!�S�x�`�H$`�: З��rA[ "៳N�APc�NX�&؜ M#w"Mk��,�,C�k3�]����(N�g�'>`2}�Ǔ�t��41����Sa{��ib�f��������ۘƜ����L*�KlTA#w�;��	�율:(ϛ����)x	f0�m�����]a�H |��	+�D��40�ћ��ڶ���Eb`0�1<mb�m��9�ٚ�s��p��xd��|�9���f~^t�Y����q�����3�M�1L*�-�Z��6��m���GT��:cTMUӿk��Q�����h�ÿ���y* )gI V)�Tx��������s# z�`uN@n ���x��?��������G���{�^ħ꾌uO���U����[���Pr ��}-ލ���=T��|���f�� ���@w�D�_��<Km�+	@�}N3̝^?�S�3��<s�0q	!̰���T��s���tx�����l���ۮ��#�P9!-N��j���j���6�Z1�[��M4,�/�ߠ���1˖�ϰ	�x��Y�1e"!��N��w90��6����P:Kc�W�al�;�H b�����e�_�B ���ܮ{\�+��v�*t����@�55	`+6š�c���+=�8g�:�/����:���/,��
����Z^ĭ���`���~ۂ�`��N�	(=�	�,)�V��X\��;0 �����\K :( ��@#^�(�벖9��N@�<���N��� �S�S�v��A��Y���H	C��h��7Ou��b�C]�*�M�0��!�5�48��|��-&Ab~�y������Z���M��g��<&��4�˝��w���X�K�3��X˩�����x��l,b��y~�s��齧Bn;�D�|��Ŕ'��S�XE�&�1����o��H��}޹�1�I5��PKIj(.2��ɍ�\c���:�;�k��8�`�YH�� iS@�Ey�@����2x�����0�֢b��؅���\h@���`�� ���~7 ��7ɧ�V ��i�O��?��O���'7�)��k{	�����ƍ��큻��w;֔݌��G�T$�h�o�P�.�C"���K�2�#wm$�[�ch���Dj�v�J Lb%`u� �qɌ�g�ʿ]���uS�HD9��2�O���C/�&1A��z<���e��7_3��O�4���͉0@I��w1��g�5$� �C��i~!Q0�!?]b�?�T��:pĜ'���>'�S�O�6N������aʈ�����M�1�1�1-US	���u
�D?/�W���M���(��)�OE���w�U�9�Z.O]:k����4f��!{�ῌ��
�g�D�k5zX���l�H "pM]��8' ��&2�T�N�����$~z�����_�sCo���������/�p����_I�z�mXS.p��#0\���b0osD�s6����
��_E �B���)�OEL;��D�o�N�#��c��T8����'��BQ��N�R;#8-� �g������8-G<N�s���1�}i+O������K���~�\�xb��l��b�}l�BML'D�D���1-c&f��	���aԧ��1c�"sMY�l�܏5������r����0o�A �����%o�t��1�G}�qr�8���	������?����Ӕ��Z����á�Ǳ��~l�I	���n��C/އ����pE`�j��Q ����Z F0�p�{, ��Ē�@M�9�t�	V.�����) ә_0s"�u�֓��&1�8|�N!+8�Ʃ�EHX�;��f :-��'����������{��6q
�x���Ӿ�y�qQ������K���^a~��t�b��4�����KTL% 1�WZ�S"R�#���$���
@���n����m.���k�-5�F�nU��H �n���`�B�]��\���\�����r�89"�b/
.)� ��{���d�:T]ׂ�Y]h�'0����X�ڎm�7��1<��u|I� �z�[ ���&�<���'���ա��?��B	�.nix����{�l�݊�%���{ ˋ�b�h7F
�W�󷢿`3z�7P ֡'gw������Z�b{6e�;��/2i��D]Q��E���	|M=-T����܏e㺿YoR��%"^ L���T�A�^�DM��Qp��tp����3�6N����n?۷��]2����x�0E'����2N&����3��B����)�:��e1e6��5�����Sa^�[���7�NDMƐ�6s1�3�4��U�� �f-Wey�G�-�s�c1+�́1V�;�OH� d_�a�?* YS
���I V��@Z����|�ꀿ �s���|q��x���t���������}�*���ৰ���-=�U��X�݃%�7b�|�p;ԥ��Н�A�D$�mK@����e�����}��2
N�N�~:8}����w�-��\3��8̠uz���\��]�N�{J zO���O�) f�'�)�5� 	�!kT��o�Z�¿=�j����e��nf�o�Ң뱢h��% �lH�,Y �
�8��pi� �&�m��5�o�W����O�՛�_�g|��ה�Wp_�wp��P�$�?������w+֔��������H��)�?z�6��ȕݹ�I	蔎���s  ٣	�SA�W�i�yO�P?�>�l����f�'��6��ό���T�'�rF����~�?��X�A�����Dr7	�Q��pX&a*&����;��0��V�	]�:��R����]�$w;��ƪ��X_z��% 3��ƼYIH�<Y�����<Ⱥ8V �/�� ���rJ�����E��4��F��At&����@@K�	;�J��N���N	�x��x������%�\��zׇ�ߝX/�Ka�w?Ƌ�`���T ���� �� �)��N��X���Z��LG b	��#��c�t�q�޳�����q���`~/��%'⏙2�_�68�>a���:=������!>�����H��rο�������f��נ�;+�w`"��_xJn�v��� ̳ ��Ld^��E�Ⱦ$Y�x��Ǟ��{I��6���@}�+�P(�k�O���e���?�Wo�<?�k<����z�5��[j������3t�����f�*=���	Pc�oS��YW���Q��j8k��)�I�Թ��{�N��~��7��C�\"�JN�3d&���mp*�l���N���8��tp �����9��L���W�Cj���t�[�����c͟ῦ�6�܎]���?���' sg[�uIܗ ��\��\R�� �iV�G����ȉ�����q�v��xa��x��Wx��Ǹ�囪O���ǰ��>l
܎u�[��K��0V|�%;ԩ  A@K@�H����Z �.f!t�p�޳�����q���>���Ɔ�����ɿ/v��3�/���)�5N�>� ��/�e����֬e*��\���Z�>�Fz61���s���`c�m���*�`E����ЕY���}q�� �K�Ậ�ˊ�s�y����r
�>�\��J) U3[P?�-� ��0?M�e״�  �kIDAT4�[����K���ߞ��G�/��+>��x��{���%�^C	�}[+��&��X[zVyaY�>Lވ%�c(�5R`�H�F��GW�Zt
�5�p�F�k���Ɲ��4�-�� �F���wƺUm�� dế]`@�
t'�.gʉs�����9�� F���y�W$��qJ��/�g��93�"�P��Y��M�.<b����[O���un0�1J��O������Z8�ϟ
��85�������s��	ⴿ	N��>߯�He���R�֏�t�a��ϰ��G{�/�j�n�ٿϳN��Gr�b<���X[vۃ�bO�㸵�x���I �8 IH�*��~��Ť�P�,���r/<�� �

��e(�J ��k*� TR �( M��$�5EH�O�D}�$�@l�/�%�o��O|q��l�O�d�\�U�{7V?��{)w`]��XM	XQ��1R�Ӓ Zb�F��Q rת�#Bw&9Jh�ZiI��" �M�'�`��y�Zz��,8���	�1�Y���A�&�,���\�D�9_"���/ju$f�~��4��>8����-���z*���s���N��	s�O��wi�:6N��g���e������9�τ�) �r��$��_�!S���@K�2�d�P�4)�{��9R�g��|_�ݏ5�-��pc�c���Y���<����O R RE .g�_Z�j�R�?� \W�  �N���ɗ�����o ��Kc���x?;���F�?�s������M_�-5�ao�c���}��ңX]rP������N��0X`I����Cw�� Z �� �% ���F �Z�s8�5p
�x��_c~���Lb���w.Lcq
ﳁS{:���Lp����i�:ט���;�0��D8}��)���3N��Bc�����g�{% j��L	9�?�V������/���lf������e�k���Oa_�q�Q�%����GZ^Ə�����9 9�ru6��(��2[ .�� �~p@}�ɘ��`AoS��_�>��k<��*�jz7�}{+î��T~+֖�J�>L߈1�(�%�0�:n@�j	X�Ntx֨kI��?� ,cЏ����
��Gpp
�x��_c~���Lb���w.Lcq
ﳁS{:���Lp����i�:ט���;�0��D8}��)���3N��Bc�����g�{% ��x�j��̥h�\�V�伿���r��D�n�,<�.����*��y��"i�:�{�o��??�`��Y�/W\��L
��aﺼX�d3��W� ����/���W�?x- �� =H��$�w8=!�����'^��#���1��.�iz	7U�<������f�)=��"E{��Аj�@[�%@Z�/��tp'��N�Z���#���)�Pt�܏e�ڿ���5(]��SR)�։2�\08X���s�y�~���.f��W����2�8-�T��ֿs�zv�������+��3���p
�S��9�����x�������9g�@/*R�������៱�������Y�w�e����/Ὼ�06�ܪZ}o�z��>��^�C�_��{����1B�>q�	�\���AȦ X�?p��׼
����4�S9 7�;	��^?�����/����ɮP���j?�=Ua{�Nl�߄5eG�B
���W0��Uu� f i	�te@� 8�� ,�H �P~/�H �8����|�����+��3���p
�S��9�����x�������9� H�翅�ߦ�%��ע׵����o�D�XŚ�ƒ۰�w���s��@�7�+���������� i�� ]��� ��� tQ "� ���c�@`� �#����|�|/'2X�����D=/��;<���o|����|�x��[���y�{7T=���۱>p3V��@A{1�����=d| Kz�/@@�
���.h�� d�ڿ�c@�S ���L�|=�}Q�-�,��w�c�`�.��p�w�G�)�O��;�u�^a���w�)�O���L&ZFL���{j���P���O������Q��'�yi��k�{]�0�ވa�&����
V�֕Q�����_�<�k�n�&���WV��-��_�_o�_ } �LBڵnd]��g�g_鵐����2�^Y���|(� _U��k��Q��f���@��>t.�P�:,�ف�ޛq(�8��:�H��m����dL>ˢ�*- N�DԄ�'��&��������������y��5��,vU݇M�wbM�f���D��yo�h�N,.�F	�16�'������ё����ђ�
͞��&�56@�[���;��G�Vd�)�qԺ0��)��of=��
�la��Z�M�SQ�p-s@���/�%B`Q�X!�W
_w �ſ�9!����{�-�����8����x!��G��<Sb
Tui�s_�Pj�#N󞊘�z�pZ��C��9��)�ߖ��e��*�֘e�I�y�C��p��3� ��	��n}k�r�߄�ϚMk�i�Q�>���14�O����/#�uS �k1���۱�h/֖���au��}�/��o��=?�[���a+!��Y@� ء�i����1f��D�vl*9��Aix�# ��ش��9��#��5>��3<��-�����j�抻�VZ(���a�D$`���c�p�6��`�֡�`-��ע-o�-BS�rE�g�B$�i8s���ξ~������&�'f �T����8Jm�����b.�)~���ۧ�)HN�C��1��{$ ���,�~���~
�B�����s���Dć���t��l�4�W���>���%h���X���o�^�.k��Ŭ���mW=�ז0������#���Y�����[��o�������NV	@"H^���58zP ������ �偑�d��7��w'�ʁ�~�g��ǻ��;Z���O����%t6�n�j�!,-ۃ����^��Ŕ����+܄�BJ �"Q��@s�2J�RE�g��;�3OK �1� p*L���; ϛ�%,4iaBi����z����ia���b.�)�f���0)(�e�~:��� �l�s���=>,`m���6��=gS ��,���~2F�y��/�/7��qK��&��������� ���Gp{5ÿ�+x��k������Yd�?yǘr�-�;�`.Q#� \�H J�C	ȣ� x��D�5Q��׉�~t��a k5�j6����Gq�x��� ��n��� Y "W��q�A��:�W<7�;|��<���l�2�=��(�;�6p+|����SFK)%;0�݆����)ڈ���,\#J�W� -" �0� u`� ��6�[�u8Z��A<�t��y�i~E:ŉ8��i~���N��
����l
�S�8��������2�g�A�6Иϟz��f�;�~:8�{�&��71����S��
�[3�8���~�^���2]��	�;�_;��
r���w2� =��J�WPk_�/- -�K���2�o7k������0���bu�al�ߎ�C�V	������/�[{ƚ?3��/9pL��m�u�� �5XDH]���U+؊���J
@���/ ֟���@�� J��O����ύ���<�����%n�4n�y �*oÚ�a���X�^����D�w+z���]lI�)J
VS�%`%%`E�t�[Z&P�ļO�⺿�� ��$>�9��VA+�d8�kZ�2x�9 �;�/3xP;�48ͯ��N�!OeFg��O���cʈ)A�f�ִ0�d�8��N��3_\�ڦ �k���R���~��1e�\�NR�1׋�����M8!���$���v(5��l��]���"��F����S�U��{����k�e����4����b�ֿ`�e��?��5��=_Ń�/��o����?f%�U���$�D h��#H  �icp��x!�G�~�VE�O� �2����?����qu�׏P��'{_���/����q��I쬽�n���QJ�a,�S�)e7`�0P��%�=�M�P��Q�TK�R�{����i��ws�]X��$�0Z �0�}�Ci�U@;�N�3y�9 �;�/�2�}Y�	gN�|�f��S���8�~*�� SFL�53h��&SaML�'@
�p*��1�)���3�+d�x78m�SP�����|�*��)�����M��i��z1�7��t�|���3`�@"8�Н
)+N�9�.k�������q�=�	�U���g��F��gM��-~�]�j�x�`0o3�
��J�!VN����C8T�9���U���"�s�/q���������J�O I��l �@���KԈ�B�\@�K����ʮ�� �"<�	5;ј҇��%p��x�vl
܄�Տ���o���y� oZV%�oi�Z��1�B@P�R-��s?����Ń=��--/b_�籭����	�CG�<pPI�x���\�����lE�w��7��h#:
7��"�Jh�_�h�[����dsVR F������y(]X_R� A�� �� "��n���wfo�,d����/�N�ZTr��MQ&�f�1!����?A�֏�`����t�Ap
2�pM����h jd������ǉ�]��=,*3e�ZTq;'�� �|Ev��0��xY�+9me��I�L֧M̶L�8`n��@�D'̐�.N�y�<~����~n��%���	?�'?�o��};���������T�Q��gYV9f�W�q�ۨ�0��X���� �Q &��Z�N�J���`?�1R����;��3���]u/ᾖo��^Ǜd��+�ԭ�'�ӡpw̼����;@��Q 2�0�Y��b
@�&�y�}� �Vs}Z+�}�OZ�x�K�R��oR~w��>3�c<��:��nm}7�?�mu�Pn��O�UGJvb� �O	��nF�-�EQ	�D`mD,� dNK �f� ��o�BE6��b���t�����69��� 6�0�͠01 n���#S`Z,Rp:q��8�c�]�f�G�Qu��iS��/�Z��2i=���1�EC�	����?�`�_��!�x��A�-N���2JNgY�@�! ����@5k�5YK���2�z;ÿ�Yԟ���;�T��/�	;���p��qG��pO�xi����Xг�''�U"�"�>�� g5Mk;6�&|��Q�������X���W��%��'�������Ow}v}G������c[�]�PA	���~��l�n�`�6�[  -�ր�g$ �00k�a����*]g���Lq*�O3h��T8�$L���� p�:!ao/�!��@��v&���)8-&���
���3��c�n�C��5x�T����/Yrj�[�BJ��Į/Y��7��q����Z�0��0����� 3X�`ND��IP*
6��M��{�Xp�D�e>O(��˦"��щt+�� X�?���k) ����-~�?�z,.��
�n�)9�����p�i�Y��S�e���'8�{��aA\R�U��`��X0c!R�q�{hP2 ���@�(��r_@��� 4G ��������_���x�-�~qǿsEK�Z�Aj��DP�䢿�x���3�?��?�����>���֪��.|3V�b¿c�0R���v(�+݊��-�%��8�
`
��
�
�9� ���|�%M�@�_�������) f�9b�!��S��9<fP�$
���a�Fτ*6+� �D�f��3�O������U[8��^����)�O���T��[���>/˩��ە���)��H�=�� u��ȉ0�\H���|�@�i��|�S�V8K`��>������8��i��	e�'ĩ�/Tfp�5u��,	�Ũ�E�{���J�{=+�[����,;�m��q8���<�i~/_�3�͊�������w�H�*���������p��zA��vX�J,a�m�޺�qo�W���7>x �F$�� VOP����q��C����ίᮮ�q��Ӹ��Al����G�,��������� " D�� - ����܏/8s��V�9=*X�k�B6�v?��pטa2�k��k��"g�� ��0�1q������|\�gsN4�y�7�����,�5f��i�hd]Wg�F�m�꧃�~t*&�\�
c_��b�v�~��7q
!�4	��"ډ0C>>�=���~�5��lfM;V $��Ϙ �6���% �H��&�	��NQD t�Gj�� 4f/A�{���J�g3��vaY�~l(�{��㶊��κ��Ž?Rc��m)䭳�Q��Թ�� �݈���hH�E[�z�W`�d3k�������|n��������:���"��!��^�r���O��G~�'�H�/��簯QN܍uU7ayhƃ���=�};1T��e��K	:��"�J *�d��M�v/�U�!��=Q�a'��:�3�z-�l6�Y|�iR��e�1`2"N8�+8�k����E��QaP)�a�k��5]+�E,�ω]�(��,b��Yoz��O�6��g�<�O����'v��Y��*.�,���{"���v�:�'B"0%@0�9fțǩ`>o��L�<�n����\l0@XC�����Yb1���w��2 ��ì���ٵm���&lC��1^�k�nƮ�#8���Y���u�K�w���k��?)��X0S��p�Ej*��=�{) ^���J�#`��*hC=�5c1zsW`ĻkC���~|��Kxf�Gx��T�Zd�J��2-% R�vBzb���]A��.�$�iÐ��l��E�C	�$l��ly����Ά������8����� �R �`�Я`�(K�`]��ǝO�M�����$Z�[�8C�he;��M�k���&#D�7},y���@|�kjXhמ6CĪ��oM-�Z�~k��֏�#�0�+�\�X���5�^bB��-M���΃ڨ&Q' �XC���Ԫ7�z�3� XZ���j�\�
�\�	@¿����a}�ǉ&#�0�M�e�S�ܞ\VY���2��l��5U\��J��0d����+=���	kL�(f��y
�Ɨ�c��|^��L! An� ���	r�Q��Qp}�y,���Z��N#A���k|΂�� vF^�ay���cy�d(n\�"r��~��r���K�r���ߓ������h?��ߊ#�O�H����߱�f��-���?3s�^.��(�.�w� e�����qy2/�"�ӌ+
9�Ⱦ�n>��R
���{u��V�?��[P�܍V���e)ڈ5�}��������.^�����Q	N��`� ��_�������^������=���`s������1�K�w�~ �j�^�@䊀��h�_��<
 ÿ9w=�=cH�0��^:�R ��O�oXĂE�
��Z�}ꀒ��U`��|O�B��NH8��ԳP0��O�zŠ#u�Qj�"ȵœ�¬��8�f�'��3A���L����8�"�&�q���2��<�+������9��n=�6'J<�ZD��NS����o��m5�����j�s~�t���SE��RD�-̚}<�j>ov�+g�k|����ؗ��hB\>M��H@����ו&�u��ڪ�W��EK��d*Xh*�OD��9�/Xraa�:X��iP���4g��Mz�{( y���h76�ބ]������m�Ʊd������2U�S�/�Jp�eE��kW���*?J�	�7���ͨM�Ds� �]*Z����Qynn�4�~��g�e�]�5b[�:5���2 ���F��?���Z��~�}������0���) �c�d'�Jv�׻=���]�]�[Б�	�y�Ж����j�L �7`!������X��F��S[XhA(�5BEf;�`���n֊zX;�}o�B��#�,�OA-n�y�B�	��+�;BuFW+���xt'�x���`T���;��p�S2�y�T�os��eR��8nS�Z����f	C�L���>�@���GIP��ZR��r0lL	0Q-Dj��F�A� 2uB�u �E��q�����Q���b��E<��m�yu���O	�����@.��:���z��s�F�>��$�y��SS���v��[Tq�F��\7Tr��2��X�S�2Vf�{l�c{���|O?�+g9�Y�N��ꢣ�Tr;�X�e��
�"巴��M��<w@���`��!�N�Y��#��<�9�\V��+JPp���Q6�
���NnGcJ?:�G1P�
��w`K�&jx�v����^� �P[�p#X�"V���H�����j��7� o�iZ:����?ឥ�`k��XWr3�U�xH� �ƈ���B_)ÿ��_�������) ( �) 2(�jfc�
@���c���3[��o^�l]����5T頕͚�4��fZ�
�x����s���g3pm�5}>ΈRǃZS#���_-p��T�S��BSÂN}��F`��1��@�u�~<2���J��6����c�pe��d*(
�0%"����w' &���=F��P���ǧFj��L�LVc}�E�G>�~����X��������^�GN��y� h�hB�� 3��1[`������	���SZ���ڲjꗚ3OX�	���T2L5UmM5�:ۢ�a_�u)T�p������f��1�ۢ�YN@����!�Բ��dR.3�P ���j��5X\���[0���y��T�|��4���%�����2=)筞 N�ǧ �Y�ϸ���3�3��������9�'�b^UF�lfs�P�Ԃ�������[�ђ�X؇k��mm���{^�Gr��緹e @Y���8��}��w�X����%;�	>>�eWw���?�����ގ�1�p(_�ѪM	n�b�f�6��|=z�֣�l�J֢˻���(^��h-X���q4卣!g>�¬�[��E usc,q{�Q�'����D�E� �> 2��ZU� �BZ5�ж�3�׏���,X�X}>%�}�z��!k��i=�S�BZP��s�C?OS�Շ:���^�5AM5YS��6�GQ��m��X�󵺌^E�H%˒	=����מ�qHof��>ڂP������n	+$���U�UP�� �~B��
��:��u�S!�g�on�>g����ԱfX'�p��d$��8��|�|�E�B���p�~�V�_�&k�EET�8m 25Q�K2��(�>����T�uh��`��>��@���s���ǎQ}]���T��WSi	�<�Ds�?�=?�����P��I�����[T ����9y�M%�����kR��F�p~R�p�E�����Oi�g�S�{($�;G����I�`�7������j�W���j���dnA�{���o���o��:�/ݸN�`e��v��=,���	9�A�w��� pj�ui���R�4@�+���W�Pz]��ը\ЈZ�F�0�%*Z��e;�=|�����^�?~������_��w�����_�??�3����~����������8f��V����"�y����WpY�$��M��������_���������������͗�	�x�x�_�����}���ДӇzw�N��Y3�dhg��<�e��(I�G��̫D��rf��֏�+}���4�����tA=�ԡla-��|,�:�/�S�$�SHmV����p�> ��ł���� sqyj=2R!O~\���p����7���gd����n�e��@��ߍ|]Ӑi#��3���.�̄���S ��4���;l���i�����\�1����g��Q�uUf���roY��5y^��X�;a�t��O��`v4�����r�&.�P�u�D�=��z�����Le��7�5�5n
�k���j%�w��6���<f��4�&��gM�	���c	
E��g-#�JJ�O�$�QZ����Q�Cd��XR���LպT�KK�{G��%�]�� ���c؟&S��-��"�E^�����L�Ձr�/>kQ(
\f�K?�� �O��7��Y��C�Cd�m'Ӑ���u#��ݔ>1��0C?
�R0��{+�^�R!R �ϖ�S��߭q
�x7	���BϪ$U����!4�-Ek�8��aе�>�3����~�/��W������^��������g�׏��?���o�Oo��w�go�o`�(* E� D[ 2/�G�%ypq��R

�,� ���!�Y��z�$�@M�Gm�/&�����F�ފ���ݟ�C/♡���W�e��W��/.�|}�/�͕����_�[�����F�|g�o񝵜
�w�c������
��x���[��o��~�7W���B�����kK��W&^�s˾�ύ}��>=�2��~�=�O5>��Uwck� V�oÒ��p���Z���G=B�4�ȕ�&�Q�D�B��J�5�i3
���$_�¢�]X(��?�D�b��-Č�����7)�o!f�I��7����c��`����T�^��̫\Ⱦ6���3��s�(�W��������SB6���>��<O�K!�(J �,
*��,��T*|�+P67d�Ϟ�爟�W�T!8�
�9�9|M3�����
f�{��z�������?�˧�w�YR~�e��"E�5Q���z��TQ4�3�#��Gȟ%oF<>.C�5G<��N��j���|2�,#�ȼ���*>�����j�ǉܙA��
!6�Wn�Bn�Bn�\�]<���5(��꩒R9u��Q�Oj��!��!��C8�o�15�kc���d��s���ɥs��I-�BM�Zb]N|����/���o�[M�P��^�}Mօ�Y79ܧd=���!��r�S{}+JԨ���Q{�ޣd�yM:_O���W"�ep�yHb�tI.�.��4�.��kyH�<�����%_]��kJ�v]y�ԙ�i��H�M8M�o��oɘk��ߖ�
����е�nVJ<Iu�YT����'7�`Q���۬�ۤ0Y���,�m��E\��B�\�B.����������eȞ����.�r+@�/s�j\�t�m<Wq߼:��k�<�(�Q��Yh�Ӊ��Q,�ل��=���+�Ǒ��p[��qW�p��p׋x��x��ex߷�T�w�w�t���D���#|~��� ��ܹs�P��We!�;S:C>���x�����͝.�;bΥ�Ȼ�,PJԊ�¹U�[Q/Wd�۵��(�ַۃ7cw�]8��0nn~w�|ww|�v|t~Um�G�_�c]/���㉞o���(O�}ӑ��_����o:�4y�������.~�L��;G���H���<���Ns_���3���;S������{�>���#��ߍ奛0\���#h�c�����P=kR5�*{%JSC�y�0$�!g��;~!2g�!�j7]����`�'�?��3�fv��g�b�����;��~.~r]�)��"�LD.xf� oN>
��p>n�%�JQ�ȇr.�/��H�\�@Ý�gJG�M��h,9�R S'���!�m*�Q5/J��
N+P���$��C2�<�Y��>�M���k��@x�?Bh���#8���)%%3b)�IY�U��Y��w6�[�b���#����n!aM�exD���0X<����(f���|����f�d]�@��dRr2��>v]�ŵ2-B֌bd�L��}n�.�3����rE�<
�|�\����zL�&r��G))KfȦ4�PҚ��QH��ڐ�V���҉�j���hSS��zlאe��k�Bf�#N�� k��J�g@i|�\.͢Z�J5ŠJQFy-��q̧����v�GY�KI��@���}��g���%ȸ�0�ӯf�_U@X�����E�5��e{D��6I��)W!�*���XȀ_xY.˃̿,�d)\����($]�F�U9X��I���(�)�y�:�i3K��eӤ�����}3m.e�ǒ��ߗ��A��@^DH�QxRj�)��y����6Tp�s�$3��_T��$�i׫L�nsV³��-�)�5���\�$�˚9���4�B�M\�-�JirY�'��5�(�.��*T�iB��n�%��7}�]۰"��/:���[���S��w?���~��8|�<�C���P�G+�����-��í���mU�F���.D �.vS <�P<��#��"�_.��,,Y˚U�B�5ImhL�A���������(ވ��]��ۏ�������Xu/��<�����p���q�\�n�����;��O;��g"�E����B�֏�"w6?�SB�ŝMQnox"�mM��֦�pK�������=�e��k��;���V�8��t}{��l�{7`�p�
Fљ?������P�]����/�B	@1���$ I�`�! �"��?3" �N! ���?� " �$�YRy���[@ٰ	��T� �bad"aT	�X��s*����&���5�!�H ?3� 	��3���m�o�q�l/�l��������{ʉOQ���Z��W��O e��T<� " S���U;�ǚ�3��emۙ
���LMܳX;��(-�Y��YE��
|	{+��l:����v
��
V��/b�^���D�ޤ��_ư����!�ӛy,�U+��y�ʬvG��Z�Tfɩ-9��9� �+�鰐SfR�L��ȥ���1����'Up=p;1�D���2�<T7��5�2��ʺΒ�,�W�k�|���eP�R�)&E��2��I?�/wJ �����?��[t]1�))��E���dkJ �-Z�d����2���$�!wE��7�w�	'r��������*��.2��${.k����\����k�\_^J�n���"��^S�Rx-%��Rv}3y�ϪG��64,�G���,�`��foƄ�e��F��ݏ�y��1�06�悛���6l-�ۊ��������n��ލ]�{,J���%�}��y�.���=p�\F	�Kug�YҌ[�����t�=�j	�]������XY�k�o��cm� ���b[�f�
݊�C�a7�1|;�P�Tށ���i՝�}���~ּ�܁U�[T����d_�m��� �[#�E�^�V��Z�͸��&��ׇcg� �o�f�����߲��6ay�z,-�NV���r9� Z<]hp���Ո��Z2��3��S�(I	���[� �[@����	@�5�p]�Fά\��
P��XI@	�CK�������~9CE`*hf!Z���"HB� a�g� T0�-�DN+�9!��&���{m���)��A'����}�Mټ25�1��p���H)[٢ �.�R��A�ß�!��"�t��Q8��g
�vmShP��5��E9R�@b�jX��?�����ߤ�|��8��i�Y�'I�E=R�\��d�?C���X�ڠ7�!B)��D���3�ߟ!���ɀ�b�2�C�_N���g�J�ہ
�I��+B��ۑ�����3���h�\�`z%EZ+���{KX.N��:��`(0��m�(���ʀ���k6%`%�5p�A6CM�53�L�1Ët�w*E ���|�*
���+r���cXx���O9�:��P �$~�"J���,�-��L�E��J�`�@|k�).On��R�Gt�[��X����x�x<e���(dR@3�"����eO!��ȴqq���{<����ʐG
f��h�%�r�p`Ns�5�P��-��#u	z2�a s���b8{#�\"[�̳�r(��cE�n�̻+s�P�bu�>���am���K T����L�^���K���O�ԅ�K܊L�H@�En���p]���yȽ�W��;#��%`^�P��)�h�@g��=c�[�N,)؀eލ��X�݁U�;��t֕]�e7`=��9�P�ߍ	�=�M�X������8��s�l|�+��-��l	��g��&�v~�v.�6.��+�YϚ�LxWb��rS<�ŅK0�?�����t�<Y�4����d�g�"�����Ϡt ��bJ Ү� 銬� ���"���B���y��稰7�_�M1��w�c�t����)H�2�WgM�H+ �[K@L+ ������Y�@J8����`���D tS�j�g��~ �	���!'~?CT�/�MFZ�욼B���0�5�|\����_�~)��D�=�Pv�m�$$m
��(�`Em'T���/d�kX�g�KS��aR͋s.�\�R�r��n���\n�\�f5��f���*EA
C.�ƚ��4�_C���)�h�P���HyV|٭���T��.�m�?���b��|**%�P���H���� ��"6!.[0�ÂH��SJ)�R�)E��2T@�)y���'�:vs�v1�<�7�m�_�l�EQ0�`0g0�% Sg������zJ��yS2�Z
�u���i?c�b?S�P�ߵ�H+@"0E@���.����q	 A�]�0�s�_�)�n�o�<�,����1�C��b�Ϥ �L�i�ʞU�)��r�������bP��l^-��F�P���P���Yԏ��!����#}	�2�Г9��,VزVb {5]k1�^G6`�k#�]�#��F=[?� - Y��M\e����t�t,��Ar�ޙ,Y`K\!�Ԍ��4���)c����Q%}9��d���5)X��Z���X�:,!�E�1Q��9��Ի��	KK,��(
Χ����d��
~�<��x=�#k'���ܻˊWbi�JL��r-�X%&_df}y2�� �s���¤��H+kͬ�4��c�W�ע"�Z���!Yƚ����V��|Z�"��i��V�9��� ���mJ@�t �'���^��c���j�����,�ʂPS:��j�c!�	�`�@���
 D<�?(?-? �M"���PF	��$�`�(gͭ��X�d#;�e�%j*�C��_��\�°�)R�"0H��c�I��*�3k��_�CW��ؑs�z9_jQ%��/�[ȗ�&|��@?Ϭ��RB$��.�M>Cޤ��_�Z�BQk���(�`m�a�)�~�q
!� �a7k���sħ��P!a�@��ib�?���($~����"�g��,����R��ʀ�S������]��d�ɺ̥L�TIz�3�n��{^,ٔ�,�p���P���)ѵŪi?Ij�"qH�k��Yk^0��.d`.�g-���9 ~�	�D`��׳9_���<���^��9_���"!��偛偋�}����'��!�e�&cß�e؏��P �z������̥<�sy
(E�o�1�]P��Vu�0B�m-�@e21�u��̤~4��3��L)h�Ak��e��	td-#�#te�Pt��� 0�3.�F���"� ����=�W0L�.E�ue��.�Z% ��Ջ�Q�ҁZ��J@S��$؞͚�k�1J�8����,E�g�s��.'+(	+0����J�p�
GF��%��L͒��db����_��Q,&C9�$�xH���]��nU�obm��CCV3�3�P�Q�j���P
k��ri.^�P!��#�k�" ���(Xx�@��gx� Ĵ���%@�PNEE�_�A���E9��B������Ѱה�)�P���g�U��L���$~ʀ�cA�E�ɚ?%@�V�R���|�j"�s_,gMZS�@���wk����v�)a��p�zI��*5c�6��Fj��A��5^iR�)Jm�P��Q�8�ɑBQ�S($�2��Ϸ�Q��e�O��b�զ ��G!k�E��f����Z(�>�)�f(j�N��(�� �T�k�t ��pr�i� ��`>��Q�àO�9_�͚���R⣜���$�3-(����w	E" D�S� H�W	�NPf�Yך�Fm"�)A̐N%)�J����� �tE���|�&" ��$1��):�� ���%���4sfү+��FI�&�t~g�3sv)�-�0��1�m�������) c�Y|]�qsޜ,/Y�Ⱥ��*9�R�c�8���"^��E��^&�C'7��mF �۔N�F�ˣur�`z�2X^1��QOh�\�r|<���	E����������tU&��si�l�]�����qa �����c� ���]����
QpM	�f�P2;�B���o�X^؀�E��Ii��u��4�14ӻh`�4�A%B[�b��0ڳ(�#��Q���@<c����mO�9��%zܣ6|L��9#d�,&C�sXx���З3�ޜ~JI��]�.G7��m�%��5�vU�o�h�Dё�g�_�d0T�V!��08���P/C��A[��yJT�?7�6{��� \����sy&\���.O,�l�
�o�b&���7����4��g�\�tQ�/MF��H��p���r�33�P@	���Kq�K�W
/m\(Y��^(M�eI�8N��ߜߦ�����ΥX�0���h&���k<���|^˚�u�����[3(3��,��䅹�s��-��e�R�
�֪�)$5�^�b���2�4�
%�B���d�*�r��̺)`�r�0)&^֪5%�]G�6��M��Ea_+���s��(|\��)`x��-($/�@��qB�|���,��l~���pY4n�9R��4�n��ǢLȡ�Rr��kC0��t��cM܁��� s;�)���p$������	�\r�����怜����LG���/�Dj�V�_$MČ�RZND���o
 q��u��lE4�Jn�t�c�Zz�'K�=�xL,�1�İub_�����IX��l��������R��$Y>���	�3�%�� ��z,���=��4.�\i�|��W!��$_������u��,���J@���� x����(|���ܬ��Y&�,�eٓ�J����5N������@'�"��D�4)�+;(ƁTnS�FI%�4n��N5�@%e���U�AȈ�j$R�a����J fϵ`�! )��K��zQ&�H���d|��I-�`I@.�*F��� �CF��}n�bA=��Q��	�ɬ!��(��Q�L!H�T4�v�������Ӛ9�-k�r@I0hg�k:�ɀ�=�5t����wfʴ�0̳�m�H������d������k����v.Ce���߂��f4�7Qd,�XS�ҡ���.�N���,e�K��;tw�����N�]��Bd��G浹H�ʍ�+����t̿$s/HRw��ws) �p&���I�����f���������d�\���+3����C	ȥ�#w%��[0ۋ�97�B1L�+n�{�+�|�F��H>���C^SCS�Z���[$����໦��Y�Ər�dJ	�@	(�i�����Y	��;�0���`c��%�e�$RH�&]�B�$���]S������4���~m%�uB��^WC��l�E6C#�<fP�Ҭ(e|McՔ��OM)����ڨM��5Bk
�=�\MAk���1��{���n.����]�� �=5eyM��|�_��],d��P���4���G���
(6	��P8QQ���.�r5ͧ�"������[\�m�X�@,	(	H����(	�"`��� k���|�� ���d�
�tJ� "����X�cD�>��d�3�|
�Fw ���:�B�H��߭I�s�Tu���r E��R�I�A��|��E,���e�ENaJGf�.}�X��ڽ����c��,�Yf͓�!��E <,sr�U�
9u��?�:B��V�,�Oy,��Xb�k|�܆62��?MZ����Ԩ��M��15"	H�0C���O�$k��HG�  -�l9p	%�2<W0T��RX�K�L��G�� kg"����0�
�UI"���d�VNۉ�tEh�4��0��4gRlZ쭙2A7���t��t��NEKFk�튶�;C]hg�k�Xض�@o�.4�@o�ސV�:�5��j��	��	��S��!5P�t~�+��x�Ԯy q�.���ܹ�șS 7k�.�����He�'_�����b�Eɘ������g	�4����0W���`���a���غ �
�ە�{���[�/�R������{O��{�$�������߳v �<`JٷU�a= �	�x�y�!3(PEJ�A�4�z�g��+�XA0�r �#�G��K%��oIkoLs��\T:mA���������{��d���`(����?bۂ�si�}uN/Yǈ@��&�����)\1���
t琢B���J�KZz��y�~�`�%��ߡC�;F�?��R]Z�Yܢ��Q�+��04M�}n�͠[�)}��.~ȂK��Vi��sM���������O��'8��1l�y]FM���-»͎�Ŏ�����t��zP��u��[��8�U���V0����}���7H�NG���ʴ��/�]`P���C�=�a��a��Lk	$@���j)S��
�>�@��#�?B�_J6ta��*o����W��v�� D�o�8��{L� �%�-��1�cB�rB�3��)�H��Ѿ�U�p[	(#I�oQR�9��M�Z����m9�@�m��/QD�c���\]#ZH �Wi��[�����c
��N]z���~Z����RFH���S֡�-H@:��J �N�1ƈ��2_����V�_ɚ G _��[2K��J^
kE)�,H@e�@ё�0�֡#]*����C��FF�[9?���B~%a�� �Z��o���	� �j��ݩ $?7萭�k��f��Xy��t
{�'� xM��&��$_��e�ש����K64����?���(��ُ�H�l����>֓�YW���aB�.�פ
�㪔�*&��2�
=���Ԇ�XZ"�h1fF�;Ux�����GG��`�L����#	=E �0��,F�=�\OI���"y$��-�YK*|y����?*���}c�O�P�R�S�a=��o�n���0tv���6��ߕ��T�z�#�lW@�d�9=7�$wB����M��� v�@�o�Ag���P�"t�9��{TT���A��(����)@��2�*�W���l�R-Z���48&���08.�o�)#�ʷ���cz�o<)� w�����g��+_� ���e��ց���S�{�A\�~.	�+B���#�����w�������_�v���p;�����y�_<n;��!�[}?�A�Q��<|��^0��rQgZ�VY���P/g]}.$��m}a[�C=��K�g�4���j�Z*PJ��K)� � ���G�;=��� HAg#�vֳD��[§c"g=�?����#�0F�F�[N{��#��64%z؀TY&7 qD���M�)
�4�N�0�j�G:��m3���G��@��[K@��WM ��:���h'շ���Sq:hZ:w��N������A�.��?�ˁۿ�����_)�!h�' :�8-9)��zQ��VU����T�GT�G���[���j� B �,s�@�ܙ��e���*�P�9ӷrCEw�@�.�	���.��������I�v��6y#/�� ����&.&����#����"6�s6�a?��?�V���n�o��oc�m��ɟ�U�X�g]Aa�(9��f��Θ�NP�G�bZ��ً��>;����zt��#  :� ,D$���*��o����VA
H@	(햙""�XP	�fB|��>����B�`�h�[�Є��# m� $�C���c����ٞFH��6Ԣ�oQ�wt�6�ٿ�#�_���OR��zW���非��H�6�Xm�U��W���P�5\l����պ�ռ���Q$|�5�����<�|��-���^��S�V��a�{����|?���q����C�a��]�B�Wye����&o����W.���or��B�W��Y�5��Nq�g�����)P.�?��4�Y�� �#�Ed�5���v��롕WRC�H@	(P%(X�˒#�r�صd�W��\J*D��$�c�����D£@��3HP�܇�����%V@(jb'-h J��j�T��Lݙ���L��1B�G6:�L	`��u%Ͼ��>W�¾��X���0k���+xc�Ĵ4�����	���"s� �o<zY�.����BZ��)I�$S�!��g�V�0����U�� ;y��*;��A�D�uxT� :�A1�!v�G�*gW24�k#��GĀ��ΟGo傝�rɎ�*�����p��Kí\���1�K�����6�u|����>���}{2b��q1�~�e腚�m�-,�yT�v�8(K}��z(JE{��"L���NFr�9*����Z�����a�;41��	տ	��Gr<u�/ !� �c#��g�K�H�$%����:�������vQ��e��bD`Z��#>*zT������[c4�-3`�Z^?�&���0C���C�N~��������C�e��m��3P��Цnv�]����]O����JxDxO���N &�V�È�>��w�K�����+����K���?�j�~�����mR��iPn�z��.�Ci�H ��v��@^��3x9��!��Ԫp=�E�T�R%�����6󭟼�?����G 4����꿑s�YhߊZ���C n���<�K6v	T�@H# ~R�1IBْ�΀׋ǯI�~�H����K���#�J��`�j<�!&]>O�e��mMB�Ihk�;�b�m��;HO	�MPH�g�������RJR����º�����Kih�Zh崟�;����)~�a�����	�@������ts��.�̗VH# ��_��J���$��� �����ɛC`$���T	(Ky�*e$��ׄA��D���!ݑ�@�)P18�H��9\��%U���C�tA`E�s�F���s�d���9��?�(�K��t^Ѱ7�o�F&��2 /�1��>�JUC�B��%�����	��n��A���'��R��d}n$��c�L���.�MG�3��S���V�lk����i�>�E ��}�P�O�$��Db�O%�k$��Z�Kf��i��		P
�@�!yD��SBJ�E@ �.�|٥�_#�	|��
T��[�����RC[�)�T�T�	 =��}�s`�mEij����m�0��S7���ۄ9�"�=$�O�?�a\��eD�o`���t����X.;=��o�w��5� l]}E�`�����>]�[�`����WJ.�������ᄾe����
 �?������Q��H��y�;��p߅J��]�D<T�
��ʾ!d�[W��"�_�M�o���M�i�W���n��k����B�������w��j�$��[ �c}��#�&�l?��'n��i�3&^K�jTϮP�T�*�2�(<�q��P0�?��ʶ ��
a)�c)���5�$���Ny�$�hI�H� Y$e���Wp�K)�M\H&~.����A��w9��	H�PH�P�rz(��h�r�=��i%�������G�L��w;���?&��6��=���?l��z�a�{����c9>=B B"�b�B�� d�����R��'�!3G��d����BJ
�i)���U�Se�0˻�#�"�BT��;������]i���yJ��3kB���P�!=��ܠ���M�\C�;���#�{ Z��J_���P����}��_�~�U���K�S闷�R�f�lg��O�'���W�`��LB��;A �}�j������;��z�ўD�H��ǟKr�T�!I/���ﴞ��F�߆�	�|&m����{�9��Jiy�Ay���ܧ�,X��De���Ud��W7��R�~�q���!a@'��H���q��@�+=¿O�R�o͸���g2�~�ꢽ�n�����C���0�r��1r=nn�w��w�
�ߣ_�z&���YhXY���_�t�����B[�)��	־���WrQ�R.kz:�7<�rI�Z���1?�u�'��&2�r�@�����_�e�7yե�G �z=�`����\S��������=�H \v��	�s��	����w��:���Se+G�d��3a�M�T��4@?�@�QK�m�R���c���vt�Ss>�3���e"v���y�
��y�4�J��K�tꕏ�@�HJ>�*��H�M y�!�w�&��T�N�АK��\�B
�)f/�J�L+9<5��槜%�]�<�R���ܕ4������)��"?)���KaL�������0% 	���\BR�~��[HJ~)%���Uf�ij6ǜ�KR��+Q�ik��"�2�@Tj*-D@;�!P?�^�*��^qhCP�����`4�D!f��C4�;����h�?��ox�o��	��i�o���� ��U�p��(n�ntp�?M�� h���W"�!G ��z�?�� ���+ ��>���xq���Ir1l �����<	��- G 4���?l���M���e���CF�_��?�� h����;3������1��v��j�2�~���v�#`-��.}WK��KP�O����-��)V 4���m%Pю�N�A=_^;G~�Ta���X�s֓�B��9�~�qU��㺆Ԑ���r��U��T�]¿��' ��`nF��K�� p[y��.��.:?�y�/2B J����s���M��&��M�:΂W��^GT�S�t��2����3������M��oɞi����o%fD@=-��!
i��v��\	� �gү}�d�  �v��H]�-�
U��ZpE�#7P��H)��� ����˥²}���S�5���߾W l�?�_ ��ʶ��;T�A�	{K+��G;�ſ� ̥%���z�$��SQ�LH�"�r�������ļUD�mPJ�U���kF�c�ӡ�_&ƝϜ��4=��+m=��t3^�t�~T���zЕ>!���@~���ڷ�?�5�M�j�_$���X�J6O�9Tw�T�@�W6�Rb= G�g�b���z��cT�J��S��	�տ	�G�&�5��>�����an��#O$��P"Ϗ$�k�y��BH�K��j��j��j��j#��M �8N��3l��[��}	����M�S��ٙ�C* ���m�#�Ǒ v���K�R���o�<�d]��G���;H��?�G�o<��z�oQ�c�6-�2բK�1���Z�Lߟ�D >[P�+� �;j��.�Cꡓ^A�R����Ͻ�>�hG��}z�ӗ߁`�\�y,7�	����m�m�,7�_ ��' �A�w�����澫�o�Kd`�� �M.���E﯆s^��Z�~�G� ?-�{��^/~E�}J(��
![f{����:��7��Yߛ�(Zrl��&�ٖ-��<�3⟒b٢�I#�)}���V.%���\Њ���̛�%�t���}H1�}��!���6�����?��s�R��I��h��&����U\*����k�;��K�����F�G�� �r�;��f-*sA��V��wif��h�?�s	�	:
K��T �R��r�j4+�ż����sBk� d��]JIf�`A2k��LK@�i	�Q	(# B_%`=��t,C
�6���4� �}NX0m��-=�NG����fg�`�^�]�H���E��M�|�HCz�tCUC��lh������&�����Y��d���6ԷRR��fR
�q8&���	��rTT�1���ܩD���T���o�_�?�ӏv�4� x��ɾ���E�s'��g��Dx?��P����J�2�V�/��{����}�>���qG:G���Da�i.�� t����:�����A�qaĎm�N�\ɽs�<G�� ��7�ػ0"�,�����v����t�i���2*s_ ���4����6�� &�~d���W�?;�ܧ�Vo�˺���+�1�g�X��0�	҅|�9�p�x�/������|]�	�An�C�m�0����w�ӹ��.w�����.//�g ��ws����`9gy�$����ߐ ���d���y�n�Gi�Y��o��:��[��\&tK	�/2���o��]ɝu�S����g��H�m[Rl�z��.[29i�:�9���H��)���`%�� �C ������� ��!?~_�W)x)���J>;&�b���YGF��+�L��r&U5�Qx� h��7y7���Dзʄ�K�m/~�F>�:a?��R�|&��g�`$`!G(e�Ԅ $�E<��A2�II/%%��6=�Ӯ�)h�h����B0���f�k�s��:hTk���*�T�:�4�	�hJ�?����jC� iB��	x=�o������i����qT���F��GC���1�w��Զ�	�By#.ŵ���"HRX҄��\�������G~r(!��G��>"�8��3�c���}�0@�ّ9��V�E$`9$�$��Ϫ��Y2�O�"��?͇���f�����`p[ ��� �> ����7y��i�7d?3- *�"/�!���D��p�}fU���/��,�?"?} |���WL�����ҩ��)Ϝs����ڄO'��@��	�A�	�a9�#a��y��(~��3�,">���k~�k~�k��M	h�� �9�z��_�
�����?���ʫ��7�۫�[n�_����1�!7��6�����r����]F]��_���Y:����x5���|�B�H qR��!����Z�#�9C۶��[f$��q���d4�}��Z�WÃ"�<��CI��CN�@� ���>�����#�I y(̠�}H�+�[�MyD ������)�%��T�*�*{���w�Ϣ�Ne¾B?�gҪP��D,�����Q�9A�}G�}H5�鿈 ,9�����Ӱ�_�*	# ��a�6� V�Lˀ+z�z��������B*�O
�����5��m�ﺝ�:',��O+&�['���Q^�9� a_�گ���Ԣ���I��ICm3q�S�W	�2U��ϯ�$���X��1��s=����@؝Z�� ��a�8���'�A@2|����+Ӈ�|� ��~�?�|h �x�H����G�C * ^ v����T��4��2`��}���>a�+}+�"食C�@z3�~(��W����{�|^d'��V��	֙�b��V��K/T�t5ͅX��JZ�kы$�(]Ġ�F��r ��k�R���C�AA[�����rY�F.k�:�[:x���!�����m�@����Ɯ�0s�?��W.��9������b��rN��4�{��G �@h" u��vSE ʹ�F J�[)�ud�!��o���Pr"Y�=� 8�����x�O Rg}����v���&n%�zΤ'�?��xd?� ���-�(�?#�?#ܙ/*��B0���-z�N�ed��T�I��	|�Q�}HZ�1�a��Ү��־�hW��G�2��4�:h���J@=�';p|� G����%����R�]d:���q����=�����?=�,,���RBr�Iɮ ��e�/V
,Ab`�-*v�T?� c��BQC�[	z��A�����4� ��}9�&�u��)[��VL��؊K��on0O���
�wy5"�ը��sT����|�@�ũ	����%��@"�%����x6]t�>g�>�E ��C�90w,	s���� +Qɮ�$���� ��6��|�P�V _�[�P�/C�Q�AtL� �T��.����N���i�z�K�9��Ԝr:�"�	k�iG/�C �	�~�F�G�GTE�J�-.���� vb#vbzyZ�"�9>]*O3�[EO��O�C0P;S�����,H�K�ڃ��r_{t}t�/s��Fv�?��'�-�[)�����-�<7�w��E`��8�c�|����)�$��򏾒F�N�ki�]JCGb<;��
���0��9��rv)�ȵ���>�6@�z���.�!p�*n�[!z��ٺ$��j?�g��z��/r���C����)p�yo��7��y\s�Uh����7A�����J�� T�ҏRG�j��*���`�wRd�ӱ��l�z)�,�i�kH��؆�Hm���^�ޒ#�-�5x-�W�T���y��H�Qw!�+�g�'�SU�i�K��6���6�g�����%���c��-���Lul���2�RQW	{?5��z�sĉPgڬ!�u�r�F��A�I��h6l��(m�y�_J��6^g[w�!��f���7���|����;--��J��B�m��Է��<�+�g�����#�Ą �� �$BE�@�@�?!�|X	Hr_jΕ � YWRH��p1�\�*�Ɂ�;�RP��2m5ZG��B ��A����5�P�^�JY{�o����*T�UC"R��FT�c�y*�*y%,�e��Q�g ����q�?� h����>D � P��.:��L�H��Ğ�p�k#�Ȇ�8P�#YW��zf��)���>E�-$`;/���e����.R��7�Ɠ 3�3m �]D`�i�#�<��$;�D�Q=$�>�0�� d���W�5�rC��" w�k�ȼC >�s�JSPm�k�[ؙ��T��������d\	p��NnL[{�a���m������iY:�h��4]�s�e`$�A��M���2#�������$�o�~v%��ԎR?H�ߦN6,�
A�tܼ�N��;o*ڙӢ�Y��V�a6�9���q��b�~��Ό�m���\w~�����-�K���j8o���r������aH��z���[���+?J�����T���i�3I��^���)|l���>��%�;�T�����֠z��^MR�u�40F�zΥ����	$J	0�	�o%��|W�X��e��/%��Rf��`���PE�k�.*�K�D��?�F��ٝ6�x��uiԾ���n|}�6�n�4��]�����ֿ�h��XZ��`C��Ol�k����_��}{L���J@⹆20aJ�Aj!*)$ ���0�\���E;ZTR>�[����E�H����9=O�p�S"ԋ�=֒�W��zB�P 8�,�\*�}e��_S�A�חC���Ϥ 9�h�I�?A��	���c��$L�o�_;��
_C~�ŶLr��=ܒ�m�>Q	ؓ��}84���@ ��,�-��!�w����XY�]�2TY��l"T6��T����棎ؑU�A���4T�E��7��%�����0DFH���h+ ;Em	�΁ÜC?�	pz�}HG�q�q���c�>��@u�W�f�b��<��L[�
��ZF"4�]&�C��u���;(m0A��o%�S�Z��ٿ�!�S�H3�V��R��I5|#����H*�C��(}�RuB���R�I��jF���S��NAo3D�i'��%���5���_��=͐*R��w��R�Z�P����?�?���G�p�����W��Ǵ~�A���=�^�V��ߩ�D@� ��OTX�e�w1�	U�+q�˿2���)|�)���iiM�7%�=�Lnu&	$ �$�M�:I}�#D�#	�Dx֓t�`�����:�P����x)��	0d�����?����◁R�eW*�
��9|�Q�?T�c�Bޝ6��
ܢ����|����wjT�.-��]����!���e��o����?a'@*�㨜h��D�r&�C&��&�#&��!�#�B���{�m/�G,	��ym�2!>��II�H��<�b�'��ܚ�x�s����3p�r�>4-6(��=��PX�R�Ǥ�t&e���r&��3��\_<��N����Q�gt��?�#���}O��i���_��U Bk�?) g��$�`y��5�����.�z�{K�H�i�#�|d��@�"1ɩ@��^\C|X?E�K)�-?����� XVYv)�"��1��N�k
���l��im	�D��z��=��ҋLu�y��"i��v%�G�9�"QY*��/�1�'_"� =�9�*�Of� �z��~�`��~�d2���&F�1��1�<��:<Ƅ�F�����W7�N����C�]�$���of?�V�Si$�I-�Z*�;)S���WR! +��*�H���FFH�Y8�F���a��sa�̈́��ޟ��v�R:�+C7w#��K~�72��[�>���rل��r�����{B�G��!|�S���|~� �E`��D @��'�;��� ,��wR/}; �y1Kx��Py��k��K�h���k��Nj`�$~Д�~C��,b{z)��8�D(	}�cD@���8�BzSH@J�ֳ�w��qz��� 
��/E���(�?��"��*P/k+�3mh�jO1Q���i4��U�� �o-u$�r�������m�����'V�������0�~:�{<�0��Ֆ D`2�@Xsc���%1�ė����{���V�4��q~Ah0�I���[�k�*9(̇M�����xbB_�߰��s;�_�C��1$���I<9���#��p�nӿ# �[ �>�$�o�G[��;�+�G{�x�/	�BI")D@�;�����S�����s�_NH��f)"^���R^I{����Y�y���2"�T���*"�Nkk%�#��I	0��kA[���a�OtP�����e� ء�͵����W�� �Y=-�9g'5*~6����2C�R�ءX�#�P�X�>=�����	�����&�c��xd�?�I�Oˁ�|ZS�	�v*
�A���O��J���i	�L��O��z�N�U��Hw��\�9�p!�ĥ�A%�L]�q-���N��9�w�w��;��K��	���˯	�w&�G�/���\���+�_+�߄����r0����*#d`��E�ߥߦ�o�$]=����T����gUYe�C�`(j/x�!=�K�J.~c������^I�.��8lLQ���'z(�N8���ȅ�f�7) ��@��T��H�K.�f&��:K>��G!=��`J��m�C�pA����`�Τ��?�5�0��]ꈾ���Lj|� l�+U����_���o��~���'���1B��H"~��1� �$����GT��"Bࢇ �?B�`��"��hS�%�M�ZE���B;@���
`ÿA�+5�B�_�ᛃ,�
PT�����8r�I� %�B�����7��G1K�uj)�MXJ	��|ң�CC{�!�Q\�: �e`�0A	�����^���&���춥� ء��O�
� �C�`gxE�+׉;��b��z�`��=��KT�T��4�D��U��T�^�2$�	�		@ ��x���Ǆ���6�N6�zp�O�zb�j����	h��f��p*ɗRK������7L	|��O�@o�^�k���H��v&��;�ԯ�`h�_&����_Ȩ񵹴�eG/#��\�t�~B_1��7��+ 0��*� �# =���D  4Xgu������
�U"@�l7�48=��#�%U�W��d#�K�+����V�mC�%�c*{]"��*�@	����J+( ���d�d��%�J	T&Zf��/�O����}�(�ս����5�]j|F��i��,6�5��2�]��O& 'r�	�t=*��D�9��i��C�'$4C ��?J��%�$$�Ǆ�K�G��&ȴY{���B�4�"�`��p1����xD��%���$��$��b��y�a=/ߌ�碽�MOz����	�,a�cZX:����_>��2��r*L�K ��V��܉d!���_h���$�I\O�#��T�QB;FxG>ށm	�ayúG��Yސ��H��-�أDm���I>;D T�%�iH���sx�%���w���=�<�B�m�RF�^ ʜCѥ0�̧��i��bF�K��%@�_[ j@m�w( � ��}�P��p�����C�]�0|e.
u��P� y��悝� W�t3�ƶ t�- ��G ���~��?h���8�쯇<t�>�7������kh�K�����	p�����ԝ/C�{�|L�����WT��"]Ģ�w��	->W3Ge�:�Q�A��y#�4d_q�k������z���p�T�z�%^�u��}��˰�oPU�w��"��_��/ZT�zEA��*���W ػ�����.v���79�q�]$��:H@	h�*��/�i�,��_��OҬ�(�����w���� �9N�)w�P�$�	�0�]H2znHD�R�z��v�sH��g]�trH1�8����s�4@�0R���k'}�T����3�B�w ���"H
�\��w�&ތA 2���u��߲�
�������3��VI��QQ+| >9��	�`t�&ӼP�O�G��O�3���E�{������� �rH� >% <�Ix"��D���lڡm��6��|7׭w���z	��~�^��[�~��b�p���*�ŐA/=��@OAf�H��G�_9�²# ��O%�nA *<��xL�{L�� @��C_{�k�}=u�)ᯧ�=�rG l5���æD?Z$� D���KH�Zz( ����4�1���A,��g���T �"( Jqs	)�'��ve)��U��`���{(@�!�׌h�ţ� ��6;K�A�ʹltT�y���9�;*��ss�s`������� �O�`�c��4��}ǿvF��}�Ì��&H�=i�?�/�U ��w�B,m��A�yL �U���4�l4��uv�A4Y��"9��6�S��"V��Y�S[־�M�+��׫��o.�k:���?�6��h����o�*}$���E��	���E�i@�uT+}K�|#U�A��[+Z�p���JX��5t�I � �]bH@T�Z�u��9�߅ OE������kI�>JZ[!f	��c�/ oQ��o��-V l�+V̙�lC�� �hM��w��]z�f	@��b1g}���_��@@�+��yq�C�y/0�X0�� D��%��m��eR �|�,�� B> ����L�K��G�1�xۈ@��x���}H�K��G�)��)"��{vf�?I�iأ�,⑟��\	�"�!`Q	�CuWr��S��]� �ӡ{ 	Ж�ȵ9����9���Ω�F���Z:�]ۃn�Z�~B`Q�\�;�1�}���Ti�	>�5�Gh����}j�O=���<���Mnid��he	l�f�iƴ�*��� ��a
�)���dG����e, >�r�\�_g�1f����^B���\��B=��L��pO�S��� ���H�k������b�Sz�I<�Z2z-}�ƾ��^{께���������g^�%��8gX졀i�0�n��� 21d! #����P	��@AC���u嬆.A�6d:ֱ=��{�����[`��|�~*l��2�j�}���GCߏ�\��S N>@ BON	z��h7�r�l���{Kd���1�����c�[:�p��	�) �>ᯧ��O	�';�6��Oů���%(�-���%�`�#�h�e[R�w�]���C@  ��Y�F�䞝�Pxz�QD
,��  ysh`��!�o	�oפ�`O��Q�@�d ó���/�K�d�����l v�#E�
H�D^I?���>y�@���zt�H��Q9�ءuى�ة贓yG���N�bF͛����H���Qi�y�Q��uюy�B��`$!C(g��=�͎֏�� (蕉��n{� 8W���O-D����F̼� �W�k�^��;��o�;s=~�.�e�/�������W�# ��1>�S�I���f	@��S-� 侒J���� ���B����(�մ���S�w��/�����M������O�D��������3[ ��;���Pt�(f�B�����vV ��ܵx��v4K ��~�,��t�O��?� ���GQ9^Kx))avҧn�����?;��㐄�L��'/�E t@�?�tЏe��t����*�^-���/�%����A	 f��(��±$�?	YB?�����_ 4�KGF r���C@���}`�E ��ᯝ��L���*qH<X�H=�p�$��m;�yt�?d�},OX~r�{z���|zH`�+� LK@		�`�Ph0��	wl 3H���A]�dxڗ��H.��\F 	�`�{a��ԭ\�!�d�Ȑ�������V��O�A��$����e�a�P�-�@��K������Pg�k�?��P)P�S��i�Ȁv���v%L�?�0	;o�2) zH��WF��(zHE�h��o�*a_�k1�2�`��`���\4�_#$`8��� ��;�O��Э�����J?H����
BUb}���"�U�|���w�j0F	� ��С|}r�G0� Ff��[I"��D������wHE��.��r��N3QD����O�m��
���2�M;ԙV-dUE����܎l��Rf��m�GD	9�SL��LV�6�-6�l�n�?W���	�C ����i�'L�s �i�D�_�wЫ�9h�!�-A�����&f`��� �[ �� ��k�G�_)@n��A
��!�1� A�'�J�ᚙ*�G���A ����" Y�i�ÞG�ɾˁ䑃� 6OC6��i	�gL@� +�V��3���oK��+}$`���*�*�9Wb�r�B�� ���t�z�^��t���m �d��ٙ�ؙt	��niSy͢�N�Rg�9�G�3�Q�Y&�O)������ց >�f��v��t��av܈O�a�ME7� mP	�Ε���aЋ-� ��� 4~���/�!����T���j߫���7�O�+��O�)# ����# ����_f��Xg&�Y�J.F�AV+e38Ї@�%�?�4!�?���C?���m!��&�@���!��%�d�����nT�
�=�7}�	G�v~�P1������t�m�����?�����o����%?������- �>�K�s�� P�?��' �� �x�A�C?����	~�<���W�0M`�+� ���N�' �|��2KT�H@��"���2ӊS��J�s<��_{�_ �@C�}- kT�)HS�g��%e�7\6	�-�=���#�Gه~~�G.�AN[���G�l#��@��+ϣN?�焿�h��P�N�" 9 � ̘ �U$`	@j�@]%�=-P;�� ��ג.�?��	���.Nrid`$#D`>�"0��� z!�����z��k�"����-�<d����W�o�O��RN��/	s��z T{cn����Rc�b��Cs�����<)`�`�۠�k�A o�@jTjU;Q�g��S�me���9�9��}!�j����:H "0,+#$���+? ?�_dT����o���w��S��?I��_/��ճ&�ߙ��M����
���P�"MQ�&�(Y7b�U#��J�0!��A�}d|���͕�> =�/�vc��	��c�K��]x�N/�q>�g�����	������4"�QPBY� �A������[���fX��65�'R2��� x��H�8cxc�M����A�̛��3~��S*�w������@=���
�'H	�	����g��C����3�>L�D�jRG��qD �(* �j�������O[��͟�$�7���X�$>��@�H-L`% �x ť ���萟'l種_�K���$ �_���z!�����h[���·��~&�W$�Ѳ$?^"�]X7����Do�r��G.�w%�|Y�c9��7���ϸ��������4�$"���B�PY�HPj��	�+�#���47+�ڪ��5��ԥ�۔2�W��Bp�5���2: p:��9mp(�йt×�\-=*�.;����.ۡbhS)t��Σ�N���1���4��6N.�zr�Q9�0���K��G�X��GAN�~�Rg�K5�J*3(^�
;�1w��C�F^R�z��C�E>�I��T�I����	�b�\���e?�~N��0@��E�9'�G��|P�Ѡ�C�W9�	o�
����<x�Ð��o���=����-�������p��x����>\����@�	n� �f8a�|�4ۣ%��H�Ag�>�8�ݘ~�D��ynB��!L�:Eh����5��3���C����"��2bZU��@[�T�J�	��6��Z�+�9���:�4��<���=��k6�E��d�~�4rD���_C N�	`���Ļ,���}�J�X�����@\���C/�c�;�$nI)�z�-��~�=�/�<ճ	�=�<�S��M����V�z1�8!<K �$� $!M�g����n�>7��˦�n���J�� 2ܗ}�g H
l~�22����-E��������T��B�RC
��9��楱V��ZQ��Q�t���ݪHw�*=����w�2@������aG�G陫�8�i�]�@�1:���C��,_������*x'��8I�h(�Á4���z�����R��Iy�/%˞C���ހy�/y�C��[��|.����Rj.*�����xX����Q�2��k
a���z��P��*U�i�@�uB[&��7�b'�}":To��D�ʯ��D�����3hR�k�F:�)�6�^�;��eX��p�y�r��㡛�ּF[Ϝ�P�kK�RC^���V�e䦄��B�!O�����S�D��a�QE{��9�Ӓ%\���B�$ۦ%�hZ���>F0���	P9�O��ZI$�O��cIS)[��C���vPb�D�R�ma��ao)#*yn7��|F��=�~���du���u�#�����_��o8��@���\���' ���U	�AL% >�<E>�T�$�G% �V�Z�������m��K�9�'�Sf�~���v�s� ���T� 	 ��
U��
��j�=Z{�N�2`%`ې~�H��6���pm18� ��X
O��ǧR|r���TB�lWŧ��3m�I*A�m�2�*���L�I�/&���ii2�Z�H{5+e-+����6���72�,� 9lWd�SE
���դ�_��AC:M���Z�9j�v.��+�CEG"���\4�ݖ4wt�4�R����*�U��R�nHq�)E�uZ�l8l�5�6���fWJ[=)m���3��K�4��3�"�f-[��|��"!P=BD��
Sm��֍*Q# �a3t#-��6�b'zk�3���#	JQ�Rq�	�v�S��SiR��f��b�[ztpK/���S.�/�/d���������_��_H+�9r��ڪaZI^J��/��J��Q"Џ	l�*�X� {x!كs1���r���:�Xy�C�i���J�%{�&�-)�ђT���Q���#~0����ix�IQ��$�CI�=���HK��ْ�. ?E���2�:�!Qud�f�С���ܾ-*	e�/p{NC���(��m��-�=�X�ҀwI�[�������8F ��c�#��	��)U�	;�S�grʎ���1zL �o�c?C,�"`�<9�]��}��9Ğ�}��?�j��Wû�V��A���Լi�v<��w%i7�gC���EG��{���>T�q�_�R�[b6�_I@��_#�	}(<\����a��>fU�<��X�	����}�����wI�%)���Lr���C��!z�@���vd)=F&�ls��g�곐�^D�>3�4�f[�q����c�^�Iw%!=��j
��S�2�[�Hwi��Jk#'�M��f��R��Pr�f^q��Ģ�Q�ƦC����;��P[w�|�vjԋ�E�JP\+K��R2�Wa�,�e���rɐc��Rᾊ�W��*�Ն�\
�M�o ��1y�!����e�ܩ�Q�JqkLi�-坎�v�R��Iu1��A_�P�M��k����:
f� i -��&v��Sm�	���}J�E/S�4�Eش	�t	�^�5r��g�KEߎ"�7<���~F0�R�_#.W�̥�.�d��I~���Jv{ }]��8�vz�=��P�R�rċ���x��^�C/'lI ���{������r/�/@�K���Y�@K��Υ���WD�vr��v�^K�ҩ�-�C�߯���S�P�@uj1�q�¼_@R>2��%}�T} )��Ͽ� �ء~t�\��xh�y��� �����S9�C8M��x������3&�d�j~����9S�GG�K�����Ӣc�{�A���#��i�'��P4���B�O�B��n0�p���d>��H}�w�������@�B�cْgyB� p)��8I��I %�+���2�O��>=�ԟ�9���Si>;���|~$-Į=w�љ?����B撂H���� ͕����aY�և1���Gͥ���\YJ��BIz�cq��NB~!㑛O{d�2�y��̋���ssy��|�#�X��ҘܲʃC�d��J�>/�{�'*Pp)�"'kU)n��ͺ��Ր
�w��ݖiQqZU:Е�P��K���FR!�t�e�T����}T�5ù�	�&���BXXZ�P�]��s�XY�����w �ۄ�Vא��Hv�-���!kh2��h�:�l#N.[Cr[m�"V��fÐ��v]�.�͚Gtk61}l�v0���D�G��#�Y�'��H��/Y�W�PU�@Y���RD��ȗ��d|2��Ȇ�$UNX���,I�ƒP��_���g��-!M�co�e�@�1�Y"�|<�$�}~�cx�����AL��]�Z�3�&{�'=�����\�zz߮D����9�� ��f?^#l�P&�-�G+>�Ň�Rx�"Em����C\2�R��7���0��K���ǈ�K�G�c�>��2�`�7W�l;5d��hL�ၙ6�v��dOZ��6��~��z/�9�X��9�H�4��B�PGjsg.!�#���G�eÂ��\�U��>ct��<�^$<���,��>�%ư�~��?.�4�{�H�q@,i����������<W1B2&;��d>���%����bNrK��2R�Ւ���V��zIjzh�oV��U�ں U�*�P�@6��C˴2��hˆ��)mw�L5^�:�� ��8bё�^�h3�H	)���t��AX���Nsk�a�JX��+uI-�|T<�+U��j�#�V�Ȭ�$��c]R�eC���@"���"�� �� �{Dd%��"�@�fg�Y�d}�7{�N T���ua��V��%�mi�+�x%����m�]C�~,K��D��EE��� �" ���iBGG;8����'$�,.gϢ@��g!��S��SB�h��-�{�C7<����y�k��QmZ��zL̏�q�V��D�򱎹O�+��Oh�h��y^��:�_�`
�	|�4??q=���%W;�9d	�<A_y�*�T�2�)�0ϴ��*��H��h��3�e ����ŏ��gP��C��Gc�<��:Rj��"P緫3m<�uٓ��ȡ�x�ቋ��~�#3�lP��ȣ�|L[[,Ϗ�#@X�͏�"+U�W*�a)-DE���,��
�"٧a�5d�Df�~��<��:��[�Sd��88����"�8� �Gc��?���\:}�3��$�8�b݌�-dL�O�V�RA�2�%("����!X�q.KJI�P%�k�uC�ய���r�Ku��Ji���U��X�RFfʒ�+#7�t��\0����'�gN-I��=��"S�DYG��"�Q�.��,+�Cl�*Q��%��8ԑ�&�S�V	��F��.�V���{�I�4�IJEʥ�D��[.��2!�4d���/�t)I����L~6>/R�a���5���[��� I3�XN�N<?�k����e���F ��6��C	����-��	��<A?w*��'�#��C������H�����ˎ���
`|�y�0ｎ���;��S"�#�k����������y��Do�����Q�^���5X����-H��D�,I�ي$��J�9���5v��)����U����#R��%�hU���I$�u���>��0W �h��
&�CO=����s�VJ�َ�fZ|��C���JϷ`��[R�S��v٥R?��L
Kc�H�A����٥S��H/�8,�HRG�t1}R<�_;#�X����?N�}<�\�;t���(,����@�c���`:�նd��4�dI)�T�'?���%5��, !ICn)�@��ICR<ǒ��{$���$f�;�1oY`ٲ�ro9&>kd��l.b8u�ȓ?��"��:]NB�ZIKxV2L3Z�y���.p[tj�0�eC����|t9YEJ���~K��W��d�
�C�E�q_��D|��Ͼ��j�Grd�l-H�����w}-GxÚ���1?�B�dyyQ���K���(�����bEV�����Y�+̯֕g��2!�aX�ϛ��Ə���}�M�o[�]����O\t�]��|��C�OaA���輻��t�c���E�>������8�-��'����������;��3}!{�����}���|�o��A��k��q/��������N�m����2�<�0��zb��-��x�=�g��:�>������Xn��`��-��`{�ރޯ����0�_��glw����輳�b�F���}�-�c�.[�۶bo�-o=^������:o�u���>��j�5��}�?�^.����gb�.�y��*��ɏ���ɺp�a�(β���k��o�΃�Z��γ���r���3��x�]v1�f��e�e�����X�&�Alp����}�����ʦaV�c�ڋmY��v���V��U3�?�t<��so�&���kms�4[<v��׹_��βA�}��ʼ�,�s��b>�]�;�/\��5�nf-o���u^k����"�:�'�    IEND�B`�   System.IO.FileInfo   OriginalPathFullPath   3C:\Users\gooey\AppData\Local\B1NARY\Saved\Slot_0.sv   3C:\Users\gooey\AppData\Local\B1NARY\Saved\Slot_0.sv   �System.Collections.Generic.Dictionary`2[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[B1NARY.Scripting.ScriptLine, B1NARY, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   VersionComparerHashSize  �System.Collections.Generic.GenericEqualityComparer`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]    	          �System.Collections.Generic.Dictionary`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   VersionComparerHashSizeKeyValuePairs  �System.Collections.Generic.GenericEqualityComparer`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]�System.Collections.Generic.KeyValuePair`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]][]   	      	   	   �System.Collections.Generic.Dictionary`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.Boolean, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   VersionComparerHashSize  �System.Collections.Generic.GenericEqualityComparer`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]    	       
   �System.Collections.Generic.Dictionary`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   VersionComparerHashSize  �System.Collections.Generic.GenericEqualityComparer`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]    	          �System.Collections.Generic.Dictionary`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.Single, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   VersionComparerHashSize  �System.Collections.Generic.GenericEqualityComparer`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]    	                jC:\Users\gooey\source\Unity\Projects\B1NARY Therin Demo Prep\Assets\StreamingAssets\Docs\PrologueStory.txt   jC:\Users\gooey\source\Unity\Projects\B1NARY Therin Demo Prep\Assets\StreamingAssets\Docs\PrologueStory.txt   �System.Collections.Generic.GenericEqualityComparer`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]       �System.Collections.Generic.GenericEqualityComparer`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]              �System.Collections.Generic.KeyValuePair`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]�����System.Collections.Generic.KeyValuePair`2[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089],[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   keyvalue   Player Name    